-- Version: 
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity MSS_025 is
	generic (
		INIT:std_logic_vector := x"0";
		ACT_UBITS:std_logic_vector := x"0";
		MEMORYFILE:string := "";
		RTC_MAIN_XTL_FREQ:real := 0.0;
		RTC_MAIN_XTL_MODE:string := "";
		DDR_CLK_FREQ:real := 0.0	);
   port( 
       CAN_RXBUS_MGPIO3A_H2F_A : out std_logic;
       CAN_RXBUS_MGPIO3A_H2F_B : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_A : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_B : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_A : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_B : out std_logic;
       CLK_CONFIG_APB : out std_logic;
       COMMS_INT : out std_logic;
       CONFIG_PRESET_N : out std_logic;
       EDAC_ERROR : out std_logic_vector(7 downto 0);
       F_FM0_RDATA : out std_logic_vector(31 downto 0);
       F_FM0_READYOUT : out std_logic;
       F_FM0_RESP : out std_logic;
       F_HM0_ADDR : out std_logic_vector(31 downto 0);
       F_HM0_ENABLE : out std_logic;
       F_HM0_SEL : out std_logic;
       F_HM0_SIZE : out std_logic_vector(1 downto 0);
       F_HM0_TRANS1 : out std_logic;
       F_HM0_WDATA : out std_logic_vector(31 downto 0);
       F_HM0_WRITE : out std_logic;
       FAB_CHRGVBUS : out std_logic;
       FAB_DISCHRGVBUS : out std_logic;
       FAB_DMPULLDOWN : out std_logic;
       FAB_DPPULLDOWN : out std_logic;
       FAB_DRVVBUS : out std_logic;
       FAB_IDPULLUP : out std_logic;
       FAB_OPMODE : out std_logic_vector(1 downto 0);
       FAB_SUSPENDM : out std_logic;
       FAB_TERMSEL : out std_logic;
       FAB_TXVALID : out std_logic;
       FAB_VCONTROL : out std_logic_vector(3 downto 0);
       FAB_VCONTROLLOADM : out std_logic;
       FAB_XCVRSEL : out std_logic_vector(1 downto 0);
       FAB_XDATAOUT : out std_logic_vector(7 downto 0);
       FACC_GLMUX_SEL : out std_logic;
       FIC32_0_MASTER : out std_logic_vector(1 downto 0);
       FIC32_1_MASTER : out std_logic_vector(1 downto 0);
       FPGA_RESET_N : out std_logic;
       GTX_CLK : out std_logic;
       H2F_INTERRUPT : out std_logic_vector(15 downto 0);
       H2F_NMI : out std_logic;
       H2FCALIB : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_A : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_B : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_A : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_B : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_A : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_B : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_A : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_B : out std_logic;
       MDCF : out std_logic;
       MDOENF : out std_logic;
       MDOF : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_A : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_B : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_A : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_B : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_A : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_B : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_A : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_B : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_A : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_B : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_A : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_B : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_A : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_B : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_A : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_B : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_A : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_B : out std_logic;
       MMUART1_DTR_MGPIO12B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_B : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_A : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_B : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_A : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_B : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_A : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_B : out std_logic;
       MPLL_LOCK : out std_logic;
       PER2_FABRIC_PADDR : out std_logic_vector(15 downto 2);
       PER2_FABRIC_PENABLE : out std_logic;
       PER2_FABRIC_PSEL : out std_logic;
       PER2_FABRIC_PWDATA : out std_logic_vector(31 downto 0);
       PER2_FABRIC_PWRITE : out std_logic;
       RTC_MATCH : out std_logic;
       SLEEPDEEP : out std_logic;
       SLEEPHOLDACK : out std_logic;
       SLEEPING : out std_logic;
       SMBALERT_NO0 : out std_logic;
       SMBALERT_NO1 : out std_logic;
       SMBSUS_NO0 : out std_logic;
       SMBSUS_NO1 : out std_logic;
       SPI0_CLK_OUT : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_A : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_B : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_A : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_B : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_A : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_B : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_A : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_B : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_A : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_B : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_A : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_B : out std_logic;
       SPI0_SS4_MGPIO19A_H2F_A : out std_logic;
       SPI0_SS5_MGPIO20A_H2F_A : out std_logic;
       SPI0_SS6_MGPIO21A_H2F_A : out std_logic;
       SPI0_SS7_MGPIO22A_H2F_A : out std_logic;
       SPI1_CLK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_A : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_B : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_A : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_B : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_A : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_B : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_A : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_B : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_A : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_B : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_A : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_B : out std_logic;
       SPI1_SS4_MGPIO17A_H2F_A : out std_logic;
       SPI1_SS5_MGPIO18A_H2F_A : out std_logic;
       SPI1_SS6_MGPIO23A_H2F_A : out std_logic;
       SPI1_SS7_MGPIO24A_H2F_A : out std_logic;
       TCGF : out std_logic_vector(9 downto 0);
       TRACECLK : out std_logic;
       TRACEDATA : out std_logic_vector(3 downto 0);
       TX_CLK : out std_logic;
       TX_ENF : out std_logic;
       TX_ERRF : out std_logic;
       TXCTL_EN_RIF : out std_logic;
       TXD_RIF : out std_logic_vector(3 downto 0);
       TXDF : out std_logic_vector(7 downto 0);
       TXEV : out std_logic;
       WDOGTIMEOUT : out std_logic;
       F_ARREADY_HREADYOUT1 : out std_logic;
       F_AWREADY_HREADYOUT0 : out std_logic;
       F_BID : out std_logic_vector(3 downto 0);
       F_BRESP_HRESP0 : out std_logic_vector(1 downto 0);
       F_BVALID : out std_logic;
       F_RDATA_HRDATA01 : out std_logic_vector(63 downto 0);
       F_RID : out std_logic_vector(3 downto 0);
       F_RLAST : out std_logic;
       F_RRESP_HRESP1 : out std_logic_vector(1 downto 0);
       F_RVALID : out std_logic;
       F_WREADY : out std_logic;
       MDDR_FABRIC_PRDATA : out std_logic_vector(15 downto 0);
       MDDR_FABRIC_PREADY : out std_logic;
       MDDR_FABRIC_PSLVERR : out std_logic;
       CAN_RXBUS_F2H_SCP : in std_logic;
       CAN_TX_EBL_F2H_SCP : in std_logic;
       CAN_TXBUS_F2H_SCP : in std_logic;
       COLF : in std_logic;
       CRSF : in std_logic;
       F2_DMAREADY : in std_logic_vector(1 downto 0);
       F2H_INTERRUPT : in std_logic_vector(15 downto 0);
       F2HCALIB : in std_logic;
       F_DMAREADY : in std_logic_vector(1 downto 0);
       F_FM0_ADDR : in std_logic_vector(31 downto 0);
       F_FM0_ENABLE : in std_logic;
       F_FM0_MASTLOCK : in std_logic;
       F_FM0_READY : in std_logic;
       F_FM0_SEL : in std_logic;
       F_FM0_SIZE : in std_logic_vector(1 downto 0);
       F_FM0_TRANS1 : in std_logic;
       F_FM0_WDATA : in std_logic_vector(31 downto 0);
       F_FM0_WRITE : in std_logic;
       F_HM0_RDATA : in std_logic_vector(31 downto 0);
       F_HM0_READY : in std_logic;
       F_HM0_RESP : in std_logic;
       FAB_AVALID : in std_logic;
       FAB_HOSTDISCON : in std_logic;
       FAB_IDDIG : in std_logic;
       FAB_LINESTATE : in std_logic_vector(1 downto 0);
       FAB_M3_RESET_N : in std_logic;
       FAB_PLL_LOCK : in std_logic;
       FAB_RXACTIVE : in std_logic;
       FAB_RXERROR : in std_logic;
       FAB_RXVALID : in std_logic;
       FAB_RXVALIDH : in std_logic;
       FAB_SESSEND : in std_logic;
       FAB_TXREADY : in std_logic;
       FAB_VBUSVALID : in std_logic;
       FAB_VSTATUS : in std_logic_vector(7 downto 0);
       FAB_XDATAIN : in std_logic_vector(7 downto 0);
       GTX_CLKPF : in std_logic;
       I2C0_BCLK : in std_logic;
       I2C0_SCL_F2H_SCP : in std_logic;
       I2C0_SDA_F2H_SCP : in std_logic;
       I2C1_BCLK : in std_logic;
       I2C1_SCL_F2H_SCP : in std_logic;
       I2C1_SDA_F2H_SCP : in std_logic;
       MDIF : in std_logic;
       MGPIO0A_F2H_GPIN : in std_logic;
       MGPIO10A_F2H_GPIN : in std_logic;
       MGPIO11A_F2H_GPIN : in std_logic;
       MGPIO11B_F2H_GPIN : in std_logic;
       MGPIO12A_F2H_GPIN : in std_logic;
       MGPIO13A_F2H_GPIN : in std_logic;
       MGPIO14A_F2H_GPIN : in std_logic;
       MGPIO15A_F2H_GPIN : in std_logic;
       MGPIO16A_F2H_GPIN : in std_logic;
       MGPIO17B_F2H_GPIN : in std_logic;
       MGPIO18B_F2H_GPIN : in std_logic;
       MGPIO19B_F2H_GPIN : in std_logic;
       MGPIO1A_F2H_GPIN : in std_logic;
       MGPIO20B_F2H_GPIN : in std_logic;
       MGPIO21B_F2H_GPIN : in std_logic;
       MGPIO22B_F2H_GPIN : in std_logic;
       MGPIO24B_F2H_GPIN : in std_logic;
       MGPIO25B_F2H_GPIN : in std_logic;
       MGPIO26B_F2H_GPIN : in std_logic;
       MGPIO27B_F2H_GPIN : in std_logic;
       MGPIO28B_F2H_GPIN : in std_logic;
       MGPIO29B_F2H_GPIN : in std_logic;
       MGPIO2A_F2H_GPIN : in std_logic;
       MGPIO30B_F2H_GPIN : in std_logic;
       MGPIO31B_F2H_GPIN : in std_logic;
       MGPIO3A_F2H_GPIN : in std_logic;
       MGPIO4A_F2H_GPIN : in std_logic;
       MGPIO5A_F2H_GPIN : in std_logic;
       MGPIO6A_F2H_GPIN : in std_logic;
       MGPIO7A_F2H_GPIN : in std_logic;
       MGPIO8A_F2H_GPIN : in std_logic;
       MGPIO9A_F2H_GPIN : in std_logic;
       MMUART0_CTS_F2H_SCP : in std_logic;
       MMUART0_DCD_F2H_SCP : in std_logic;
       MMUART0_DSR_F2H_SCP : in std_logic;
       MMUART0_DTR_F2H_SCP : in std_logic;
       MMUART0_RI_F2H_SCP : in std_logic;
       MMUART0_RTS_F2H_SCP : in std_logic;
       MMUART0_RXD_F2H_SCP : in std_logic;
       MMUART0_SCK_F2H_SCP : in std_logic;
       MMUART0_TXD_F2H_SCP : in std_logic;
       MMUART1_CTS_F2H_SCP : in std_logic;
       MMUART1_DCD_F2H_SCP : in std_logic;
       MMUART1_DSR_F2H_SCP : in std_logic;
       MMUART1_RI_F2H_SCP : in std_logic;
       MMUART1_RTS_F2H_SCP : in std_logic;
       MMUART1_RXD_F2H_SCP : in std_logic;
       MMUART1_SCK_F2H_SCP : in std_logic;
       MMUART1_TXD_F2H_SCP : in std_logic;
       PER2_FABRIC_PRDATA : in std_logic_vector(31 downto 0);
       PER2_FABRIC_PREADY : in std_logic;
       PER2_FABRIC_PSLVERR : in std_logic;
       RCGF : in std_logic_vector(9 downto 0);
       RX_CLKPF : in std_logic;
       RX_DVF : in std_logic;
       RX_ERRF : in std_logic;
       RX_EV : in std_logic;
       RXDF : in std_logic_vector(7 downto 0);
       SLEEPHOLDREQ : in std_logic;
       SMBALERT_NI0 : in std_logic;
       SMBALERT_NI1 : in std_logic;
       SMBSUS_NI0 : in std_logic;
       SMBSUS_NI1 : in std_logic;
       SPI0_CLK_IN : in std_logic;
       SPI0_SDI_F2H_SCP : in std_logic;
       SPI0_SDO_F2H_SCP : in std_logic;
       SPI0_SS0_F2H_SCP : in std_logic;
       SPI0_SS1_F2H_SCP : in std_logic;
       SPI0_SS2_F2H_SCP : in std_logic;
       SPI0_SS3_F2H_SCP : in std_logic;
       SPI1_CLK_IN : in std_logic;
       SPI1_SDI_F2H_SCP : in std_logic;
       SPI1_SDO_F2H_SCP : in std_logic;
       SPI1_SS0_F2H_SCP : in std_logic;
       SPI1_SS1_F2H_SCP : in std_logic;
       SPI1_SS2_F2H_SCP : in std_logic;
       SPI1_SS3_F2H_SCP : in std_logic;
       TX_CLKPF : in std_logic;
       USER_MSS_GPIO_RESET_N : in std_logic;
       USER_MSS_RESET_N : in std_logic;
       XCLK_FAB : in std_logic;
       CLK_BASE : in std_logic;
       CLK_MDDR_APB : in std_logic;
       F_ARADDR_HADDR1 : in std_logic_vector(31 downto 0);
       F_ARBURST_HTRANS1 : in std_logic_vector(1 downto 0);
       F_ARID_HSEL1 : in std_logic_vector(3 downto 0);
       F_ARLEN_HBURST1 : in std_logic_vector(3 downto 0);
       F_ARLOCK_HMASTLOCK1 : in std_logic_vector(1 downto 0);
       F_ARSIZE_HSIZE1 : in std_logic_vector(1 downto 0);
       F_ARVALID_HWRITE1 : in std_logic;
       F_AWADDR_HADDR0 : in std_logic_vector(31 downto 0);
       F_AWBURST_HTRANS0 : in std_logic_vector(1 downto 0);
       F_AWID_HSEL0 : in std_logic_vector(3 downto 0);
       F_AWLEN_HBURST0 : in std_logic_vector(3 downto 0);
       F_AWLOCK_HMASTLOCK0 : in std_logic_vector(1 downto 0);
       F_AWSIZE_HSIZE0 : in std_logic_vector(1 downto 0);
       F_AWVALID_HWRITE0 : in std_logic;
       F_BREADY : in std_logic;
       F_RMW_AXI : in std_logic;
       F_RREADY : in std_logic;
       F_WDATA_HWDATA01 : in std_logic_vector(63 downto 0);
       F_WID_HREADY01 : in std_logic_vector(3 downto 0);
       F_WLAST : in std_logic;
       F_WSTRB : in std_logic_vector(7 downto 0);
       F_WVALID : in std_logic;
       FPGA_MDDR_ARESET_N : in std_logic;
       MDDR_FABRIC_PADDR : in std_logic_vector(10 downto 2);
       MDDR_FABRIC_PENABLE : in std_logic;
       MDDR_FABRIC_PSEL : in std_logic;
       MDDR_FABRIC_PWDATA : in std_logic_vector(15 downto 0);
       MDDR_FABRIC_PWRITE : in std_logic;
       PRESET_N : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN : in std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN : in std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN : in std_logic;
       DM_IN : in std_logic_vector(2 downto 0);
       DRAM_DQ_IN : in std_logic_vector(17 downto 0);
       DRAM_DQS_IN : in std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_IN : in std_logic_vector(1 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN : in std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN : in std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN : in std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN : in std_logic;
       MGPIO25A_IN : in std_logic;
       MGPIO26A_IN : in std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN : in std_logic;
       MMUART0_DCD_MGPIO22B_IN : in std_logic;
       MMUART0_DSR_MGPIO20B_IN : in std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN : in std_logic;
       MMUART0_RI_MGPIO21B_IN : in std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN : in std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_IN : in std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN : in std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN : in std_logic;
       MMUART1_CTS_MGPIO13B_IN : in std_logic;
       MMUART1_DCD_MGPIO16B_IN : in std_logic;
       MMUART1_DSR_MGPIO14B_IN : in std_logic;
       MMUART1_DTR_MGPIO12B_IN : in std_logic;
       MMUART1_RI_MGPIO15B_IN : in std_logic;
       MMUART1_RTS_MGPIO11B_IN : in std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN : in std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN : in std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN : in std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN : in std_logic;
       RGMII_MDC_RMII_MDC_IN : in std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN : in std_logic;
       RGMII_RX_CLK_IN : in std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN : in std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN : in std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN : in std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN : in std_logic;
       RGMII_RXD3_USBB_DATA4_IN : in std_logic;
       RGMII_TX_CLK_IN : in std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN : in std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN : in std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN : in std_logic;
       RGMII_TXD2_USBB_DATA5_IN : in std_logic;
       RGMII_TXD3_USBB_DATA6_IN : in std_logic;
       SPI0_SCK_USBA_XCLK_IN : in std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_IN : in std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_IN : in std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_IN : in std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN : in std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN : in std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN : in std_logic;
       SPI0_SS4_MGPIO19A_IN : in std_logic;
       SPI0_SS5_MGPIO20A_IN : in std_logic;
       SPI0_SS6_MGPIO21A_IN : in std_logic;
       SPI0_SS7_MGPIO22A_IN : in std_logic;
       SPI1_SCK_IN : in std_logic;
       SPI1_SDI_MGPIO11A_IN : in std_logic;
       SPI1_SDO_MGPIO12A_IN : in std_logic;
       SPI1_SS0_MGPIO13A_IN : in std_logic;
       SPI1_SS1_MGPIO14A_IN : in std_logic;
       SPI1_SS2_MGPIO15A_IN : in std_logic;
       SPI1_SS3_MGPIO16A_IN : in std_logic;
       SPI1_SS4_MGPIO17A_IN : in std_logic;
       SPI1_SS5_MGPIO18A_IN : in std_logic;
       SPI1_SS6_MGPIO23A_IN : in std_logic;
       SPI1_SS7_MGPIO24A_IN : in std_logic;
       USBC_XCLK_IN : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT : out std_logic;
       DRAM_ADDR : out std_logic_vector(15 downto 0);
       DRAM_BA : out std_logic_vector(2 downto 0);
       DRAM_CASN : out std_logic;
       DRAM_CKE : out std_logic;
       DRAM_CLK : out std_logic;
       DRAM_CSN : out std_logic;
       DRAM_DM_RDQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_DQ_OUT : out std_logic_vector(17 downto 0);
       DRAM_DQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_OUT : out std_logic_vector(1 downto 0);
       DRAM_ODT : out std_logic;
       DRAM_RASN : out std_logic;
       DRAM_RSTN : out std_logic;
       DRAM_WEN : out std_logic;
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT : out std_logic;
       MGPIO25A_OUT : out std_logic;
       MGPIO26A_OUT : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT : out std_logic;
       MMUART0_DCD_MGPIO22B_OUT : out std_logic;
       MMUART0_DSR_MGPIO20B_OUT : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT : out std_logic;
       MMUART0_RI_MGPIO21B_OUT : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT : out std_logic;
       MMUART1_CTS_MGPIO13B_OUT : out std_logic;
       MMUART1_DCD_MGPIO16B_OUT : out std_logic;
       MMUART1_DSR_MGPIO14B_OUT : out std_logic;
       MMUART1_DTR_MGPIO12B_OUT : out std_logic;
       MMUART1_RI_MGPIO15B_OUT : out std_logic;
       MMUART1_RTS_MGPIO11B_OUT : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT : out std_logic;
       RGMII_MDC_RMII_MDC_OUT : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT : out std_logic;
       RGMII_RX_CLK_OUT : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT : out std_logic;
       RGMII_RXD3_USBB_DATA4_OUT : out std_logic;
       RGMII_TX_CLK_OUT : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT : out std_logic;
       RGMII_TXD2_USBB_DATA5_OUT : out std_logic;
       RGMII_TXD3_USBB_DATA6_OUT : out std_logic;
       SPI0_SCK_USBA_XCLK_OUT : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OUT : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT : out std_logic;
       SPI0_SS4_MGPIO19A_OUT : out std_logic;
       SPI0_SS5_MGPIO20A_OUT : out std_logic;
       SPI0_SS6_MGPIO21A_OUT : out std_logic;
       SPI0_SS7_MGPIO22A_OUT : out std_logic;
       SPI1_SCK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_OUT : out std_logic;
       SPI1_SDO_MGPIO12A_OUT : out std_logic;
       SPI1_SS0_MGPIO13A_OUT : out std_logic;
       SPI1_SS1_MGPIO14A_OUT : out std_logic;
       SPI1_SS2_MGPIO15A_OUT : out std_logic;
       SPI1_SS3_MGPIO16A_OUT : out std_logic;
       SPI1_SS4_MGPIO17A_OUT : out std_logic;
       SPI1_SS5_MGPIO18A_OUT : out std_logic;
       SPI1_SS6_MGPIO23A_OUT : out std_logic;
       SPI1_SS7_MGPIO24A_OUT : out std_logic;
       USBC_XCLK_OUT : out std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE : out std_logic;
       DM_OE : out std_logic_vector(2 downto 0);
       DRAM_DQ_OE : out std_logic_vector(17 downto 0);
       DRAM_DQS_OE : out std_logic_vector(2 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE : out std_logic;
       MGPIO25A_OE : out std_logic;
       MGPIO26A_OE : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE : out std_logic;
       MMUART0_DCD_MGPIO22B_OE : out std_logic;
       MMUART0_DSR_MGPIO20B_OE : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE : out std_logic;
       MMUART0_RI_MGPIO21B_OE : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OE : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE : out std_logic;
       MMUART1_CTS_MGPIO13B_OE : out std_logic;
       MMUART1_DCD_MGPIO16B_OE : out std_logic;
       MMUART1_DSR_MGPIO14B_OE : out std_logic;
       MMUART1_DTR_MGPIO12B_OE : out std_logic;
       MMUART1_RI_MGPIO15B_OE : out std_logic;
       MMUART1_RTS_MGPIO11B_OE : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE : out std_logic;
       RGMII_MDC_RMII_MDC_OE : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE : out std_logic;
       RGMII_RX_CLK_OE : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE : out std_logic;
       RGMII_RXD3_USBB_DATA4_OE : out std_logic;
       RGMII_TX_CLK_OE : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE : out std_logic;
       RGMII_TXD2_USBB_DATA5_OE : out std_logic;
       RGMII_TXD3_USBB_DATA6_OE : out std_logic;
       SPI0_SCK_USBA_XCLK_OE : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OE : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OE : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OE : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE : out std_logic;
       SPI0_SS4_MGPIO19A_OE : out std_logic;
       SPI0_SS5_MGPIO20A_OE : out std_logic;
       SPI0_SS6_MGPIO21A_OE : out std_logic;
       SPI0_SS7_MGPIO22A_OE : out std_logic;
       SPI1_SCK_OE : out std_logic;
       SPI1_SDI_MGPIO11A_OE : out std_logic;
       SPI1_SDO_MGPIO12A_OE : out std_logic;
       SPI1_SS0_MGPIO13A_OE : out std_logic;
       SPI1_SS1_MGPIO14A_OE : out std_logic;
       SPI1_SS2_MGPIO15A_OE : out std_logic;
       SPI1_SS3_MGPIO16A_OE : out std_logic;
       SPI1_SS4_MGPIO17A_OE : out std_logic;
       SPI1_SS5_MGPIO18A_OE : out std_logic;
       SPI1_SS6_MGPIO23A_OE : out std_logic;
       SPI1_SS7_MGPIO24A_OE : out std_logic;
       USBC_XCLK_OE : out std_logic
   );
end MSS_025;
architecture DEF_ARCH of MSS_025 is 

   attribute syn_black_box : boolean;
   attribute syn_black_box of DEF_ARCH : architecture is true;
   attribute syn_tsu0: string;
   attribute syn_tsu0 of DEF_ARCH : architecture is " F2HCALIB->CLK_BASE = 1.331";
   attribute syn_tsu1: string;
   attribute syn_tsu1 of DEF_ARCH : architecture is " F2H_INTERRUPT[0]->CLK_BASE = 0.971";
   attribute syn_tsu2: string;
   attribute syn_tsu2 of DEF_ARCH : architecture is " F2H_INTERRUPT[10]->CLK_BASE = 1.103";
   attribute syn_tsu3: string;
   attribute syn_tsu3 of DEF_ARCH : architecture is " F2H_INTERRUPT[11]->CLK_BASE = 1.038";
   attribute syn_tsu4: string;
   attribute syn_tsu4 of DEF_ARCH : architecture is " F2H_INTERRUPT[12]->CLK_BASE = 1.024";
   attribute syn_tsu5: string;
   attribute syn_tsu5 of DEF_ARCH : architecture is " F2H_INTERRUPT[13]->CLK_BASE = 1.007";
   attribute syn_tsu6: string;
   attribute syn_tsu6 of DEF_ARCH : architecture is " F2H_INTERRUPT[14]->CLK_BASE = 1.037";
   attribute syn_tsu7: string;
   attribute syn_tsu7 of DEF_ARCH : architecture is " F2H_INTERRUPT[15]->CLK_BASE = 1.009";
   attribute syn_tsu8: string;
   attribute syn_tsu8 of DEF_ARCH : architecture is " F2H_INTERRUPT[1]->CLK_BASE = 0.978";
   attribute syn_tsu9: string;
   attribute syn_tsu9 of DEF_ARCH : architecture is " F2H_INTERRUPT[2]->CLK_BASE = 1.04";
   attribute syn_tsu10: string;
   attribute syn_tsu10 of DEF_ARCH : architecture is " F2H_INTERRUPT[3]->CLK_BASE = 0.972";
   attribute syn_tsu11: string;
   attribute syn_tsu11 of DEF_ARCH : architecture is " F2H_INTERRUPT[4]->CLK_BASE = 1.019";
   attribute syn_tsu12: string;
   attribute syn_tsu12 of DEF_ARCH : architecture is " F2H_INTERRUPT[5]->CLK_BASE = 1.06";
   attribute syn_tsu13: string;
   attribute syn_tsu13 of DEF_ARCH : architecture is " F2H_INTERRUPT[6]->CLK_BASE = 1.01";
   attribute syn_tsu14: string;
   attribute syn_tsu14 of DEF_ARCH : architecture is " F2H_INTERRUPT[7]->CLK_BASE = 1.005";
   attribute syn_tsu15: string;
   attribute syn_tsu15 of DEF_ARCH : architecture is " F2H_INTERRUPT[8]->CLK_BASE = 1.042";
   attribute syn_tsu16: string;
   attribute syn_tsu16 of DEF_ARCH : architecture is " F2H_INTERRUPT[9]->CLK_BASE = 0.995";
   attribute syn_tsu17: string;
   attribute syn_tsu17 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[0]->CLK_BASE = 1.53";
   attribute syn_tsu18: string;
   attribute syn_tsu18 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[10]->CLK_BASE = 1.63";
   attribute syn_tsu19: string;
   attribute syn_tsu19 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[11]->CLK_BASE = 1.482";
   attribute syn_tsu20: string;
   attribute syn_tsu20 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[12]->CLK_BASE = 1.5";
   attribute syn_tsu21: string;
   attribute syn_tsu21 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[13]->CLK_BASE = 1.566";
   attribute syn_tsu22: string;
   attribute syn_tsu22 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[14]->CLK_BASE = 1.492";
   attribute syn_tsu23: string;
   attribute syn_tsu23 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[15]->CLK_BASE = 1.513";
   attribute syn_tsu24: string;
   attribute syn_tsu24 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[16]->CLK_BASE = 1.664";
   attribute syn_tsu25: string;
   attribute syn_tsu25 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[17]->CLK_BASE = 1.567";
   attribute syn_tsu26: string;
   attribute syn_tsu26 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[18]->CLK_BASE = 1.651";
   attribute syn_tsu27: string;
   attribute syn_tsu27 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[19]->CLK_BASE = 1.68";
   attribute syn_tsu28: string;
   attribute syn_tsu28 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[1]->CLK_BASE = 1.398";
   attribute syn_tsu29: string;
   attribute syn_tsu29 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[20]->CLK_BASE = 1.663";
   attribute syn_tsu30: string;
   attribute syn_tsu30 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[21]->CLK_BASE = 1.591";
   attribute syn_tsu31: string;
   attribute syn_tsu31 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[22]->CLK_BASE = 1.598";
   attribute syn_tsu32: string;
   attribute syn_tsu32 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[23]->CLK_BASE = 1.675";
   attribute syn_tsu33: string;
   attribute syn_tsu33 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[24]->CLK_BASE = 1.569";
   attribute syn_tsu34: string;
   attribute syn_tsu34 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[25]->CLK_BASE = 1.653";
   attribute syn_tsu35: string;
   attribute syn_tsu35 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[26]->CLK_BASE = 1.633";
   attribute syn_tsu36: string;
   attribute syn_tsu36 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[27]->CLK_BASE = 1.633";
   attribute syn_tsu37: string;
   attribute syn_tsu37 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[28]->CLK_BASE = 1.604";
   attribute syn_tsu38: string;
   attribute syn_tsu38 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[29]->CLK_BASE = 1.675";
   attribute syn_tsu39: string;
   attribute syn_tsu39 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[2]->CLK_BASE = 1.53";
   attribute syn_tsu40: string;
   attribute syn_tsu40 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[30]->CLK_BASE = 1.574";
   attribute syn_tsu41: string;
   attribute syn_tsu41 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[31]->CLK_BASE = 1.522";
   attribute syn_tsu42: string;
   attribute syn_tsu42 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[3]->CLK_BASE = 1.56";
   attribute syn_tsu43: string;
   attribute syn_tsu43 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[4]->CLK_BASE = 1.717";
   attribute syn_tsu44: string;
   attribute syn_tsu44 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[5]->CLK_BASE = 1.546";
   attribute syn_tsu45: string;
   attribute syn_tsu45 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[6]->CLK_BASE = 1.513";
   attribute syn_tsu46: string;
   attribute syn_tsu46 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[7]->CLK_BASE = 1.543";
   attribute syn_tsu47: string;
   attribute syn_tsu47 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[8]->CLK_BASE = 1.624";
   attribute syn_tsu48: string;
   attribute syn_tsu48 of DEF_ARCH : architecture is " F_ARADDR_HADDR1[9]->CLK_BASE = 1.567";
   attribute syn_tsu49: string;
   attribute syn_tsu49 of DEF_ARCH : architecture is " F_ARBURST_HTRANS1[1]->CLK_BASE = 1.646";
   attribute syn_tsu50: string;
   attribute syn_tsu50 of DEF_ARCH : architecture is " F_ARID_HSEL1[0]->CLK_BASE = 1.636";
   attribute syn_tsu51: string;
   attribute syn_tsu51 of DEF_ARCH : architecture is " F_ARLOCK_HMASTLOCK1[0]->CLK_BASE = 1.605";
   attribute syn_tsu52: string;
   attribute syn_tsu52 of DEF_ARCH : architecture is " F_ARSIZE_HSIZE1[0]->CLK_BASE = 1.018";
   attribute syn_tsu53: string;
   attribute syn_tsu53 of DEF_ARCH : architecture is " F_ARSIZE_HSIZE1[1]->CLK_BASE = 1.434";
   attribute syn_tsu54: string;
   attribute syn_tsu54 of DEF_ARCH : architecture is " F_ARVALID_HWRITE1->CLK_BASE = 1.72";
   attribute syn_tsu55: string;
   attribute syn_tsu55 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[0]->CLK_BASE = 1.535";
   attribute syn_tsu56: string;
   attribute syn_tsu56 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[10]->CLK_BASE = 1.695";
   attribute syn_tsu57: string;
   attribute syn_tsu57 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[11]->CLK_BASE = 1.739";
   attribute syn_tsu58: string;
   attribute syn_tsu58 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[12]->CLK_BASE = 1.651";
   attribute syn_tsu59: string;
   attribute syn_tsu59 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[13]->CLK_BASE = 1.657";
   attribute syn_tsu60: string;
   attribute syn_tsu60 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[14]->CLK_BASE = 1.682";
   attribute syn_tsu61: string;
   attribute syn_tsu61 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[15]->CLK_BASE = 1.654";
   attribute syn_tsu62: string;
   attribute syn_tsu62 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[16]->CLK_BASE = 1.683";
   attribute syn_tsu63: string;
   attribute syn_tsu63 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[17]->CLK_BASE = 1.699";
   attribute syn_tsu64: string;
   attribute syn_tsu64 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[18]->CLK_BASE = 1.682";
   attribute syn_tsu65: string;
   attribute syn_tsu65 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[19]->CLK_BASE = 1.65";
   attribute syn_tsu66: string;
   attribute syn_tsu66 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[1]->CLK_BASE = 1.57";
   attribute syn_tsu67: string;
   attribute syn_tsu67 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[20]->CLK_BASE = 1.64";
   attribute syn_tsu68: string;
   attribute syn_tsu68 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[21]->CLK_BASE = 1.711";
   attribute syn_tsu69: string;
   attribute syn_tsu69 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[22]->CLK_BASE = 1.601";
   attribute syn_tsu70: string;
   attribute syn_tsu70 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[23]->CLK_BASE = 1.576";
   attribute syn_tsu71: string;
   attribute syn_tsu71 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[24]->CLK_BASE = 1.653";
   attribute syn_tsu72: string;
   attribute syn_tsu72 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[25]->CLK_BASE = 1.68";
   attribute syn_tsu73: string;
   attribute syn_tsu73 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[26]->CLK_BASE = 1.578";
   attribute syn_tsu74: string;
   attribute syn_tsu74 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[27]->CLK_BASE = 1.603";
   attribute syn_tsu75: string;
   attribute syn_tsu75 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[28]->CLK_BASE = 1.606";
   attribute syn_tsu76: string;
   attribute syn_tsu76 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[29]->CLK_BASE = 1.608";
   attribute syn_tsu77: string;
   attribute syn_tsu77 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[2]->CLK_BASE = 1.534";
   attribute syn_tsu78: string;
   attribute syn_tsu78 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[30]->CLK_BASE = 1.606";
   attribute syn_tsu79: string;
   attribute syn_tsu79 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[31]->CLK_BASE = 1.65";
   attribute syn_tsu80: string;
   attribute syn_tsu80 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[3]->CLK_BASE = 1.468";
   attribute syn_tsu81: string;
   attribute syn_tsu81 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[4]->CLK_BASE = 1.636";
   attribute syn_tsu82: string;
   attribute syn_tsu82 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[5]->CLK_BASE = 1.614";
   attribute syn_tsu83: string;
   attribute syn_tsu83 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[6]->CLK_BASE = 1.609";
   attribute syn_tsu84: string;
   attribute syn_tsu84 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[7]->CLK_BASE = 1.589";
   attribute syn_tsu85: string;
   attribute syn_tsu85 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[8]->CLK_BASE = 1.625";
   attribute syn_tsu86: string;
   attribute syn_tsu86 of DEF_ARCH : architecture is " F_AWADDR_HADDR0[9]->CLK_BASE = 1.661";
   attribute syn_tsu87: string;
   attribute syn_tsu87 of DEF_ARCH : architecture is " F_AWBURST_HTRANS0[1]->CLK_BASE = 1.696";
   attribute syn_tsu88: string;
   attribute syn_tsu88 of DEF_ARCH : architecture is " F_AWID_HSEL0[0]->CLK_BASE = 1.731";
   attribute syn_tsu89: string;
   attribute syn_tsu89 of DEF_ARCH : architecture is " F_AWLOCK_HMASTLOCK0[0]->CLK_BASE = 1.728";
   attribute syn_tsu90: string;
   attribute syn_tsu90 of DEF_ARCH : architecture is " F_AWSIZE_HSIZE0[0]->CLK_BASE = 1.204";
   attribute syn_tsu91: string;
   attribute syn_tsu91 of DEF_ARCH : architecture is " F_AWSIZE_HSIZE0[1]->CLK_BASE = 1.374";
   attribute syn_tsu92: string;
   attribute syn_tsu92 of DEF_ARCH : architecture is " F_AWVALID_HWRITE0->CLK_BASE = 1.68";
   attribute syn_tsu93: string;
   attribute syn_tsu93 of DEF_ARCH : architecture is " F_FM0_ADDR[0]->CLK_BASE = 0.976";
   attribute syn_tsu94: string;
   attribute syn_tsu94 of DEF_ARCH : architecture is " F_FM0_ADDR[10]->CLK_BASE = 1.007";
   attribute syn_tsu95: string;
   attribute syn_tsu95 of DEF_ARCH : architecture is " F_FM0_ADDR[11]->CLK_BASE = 1.031";
   attribute syn_tsu96: string;
   attribute syn_tsu96 of DEF_ARCH : architecture is " F_FM0_ADDR[12]->CLK_BASE = 1.063";
   attribute syn_tsu97: string;
   attribute syn_tsu97 of DEF_ARCH : architecture is " F_FM0_ADDR[13]->CLK_BASE = 1.161";
   attribute syn_tsu98: string;
   attribute syn_tsu98 of DEF_ARCH : architecture is " F_FM0_ADDR[14]->CLK_BASE = 1.044";
   attribute syn_tsu99: string;
   attribute syn_tsu99 of DEF_ARCH : architecture is " F_FM0_ADDR[15]->CLK_BASE = 1.16";
   attribute syn_tsu100: string;
   attribute syn_tsu100 of DEF_ARCH : architecture is " F_FM0_ADDR[16]->CLK_BASE = 1.033";
   attribute syn_tsu101: string;
   attribute syn_tsu101 of DEF_ARCH : architecture is " F_FM0_ADDR[17]->CLK_BASE = 0.6";
   attribute syn_tsu102: string;
   attribute syn_tsu102 of DEF_ARCH : architecture is " F_FM0_ADDR[18]->CLK_BASE = 0.791";
   attribute syn_tsu103: string;
   attribute syn_tsu103 of DEF_ARCH : architecture is " F_FM0_ADDR[19]->CLK_BASE = 0.573";
   attribute syn_tsu104: string;
   attribute syn_tsu104 of DEF_ARCH : architecture is " F_FM0_ADDR[1]->CLK_BASE = 0.998";
   attribute syn_tsu105: string;
   attribute syn_tsu105 of DEF_ARCH : architecture is " F_FM0_ADDR[20]->CLK_BASE = 0.595";
   attribute syn_tsu106: string;
   attribute syn_tsu106 of DEF_ARCH : architecture is " F_FM0_ADDR[21]->CLK_BASE = 0.546";
   attribute syn_tsu107: string;
   attribute syn_tsu107 of DEF_ARCH : architecture is " F_FM0_ADDR[22]->CLK_BASE = 0.592";
   attribute syn_tsu108: string;
   attribute syn_tsu108 of DEF_ARCH : architecture is " F_FM0_ADDR[23]->CLK_BASE = 0.608";
   attribute syn_tsu109: string;
   attribute syn_tsu109 of DEF_ARCH : architecture is " F_FM0_ADDR[24]->CLK_BASE = 0.601";
   attribute syn_tsu110: string;
   attribute syn_tsu110 of DEF_ARCH : architecture is " F_FM0_ADDR[25]->CLK_BASE = 0.692";
   attribute syn_tsu111: string;
   attribute syn_tsu111 of DEF_ARCH : architecture is " F_FM0_ADDR[26]->CLK_BASE = 0.735";
   attribute syn_tsu112: string;
   attribute syn_tsu112 of DEF_ARCH : architecture is " F_FM0_ADDR[27]->CLK_BASE = 0.749";
   attribute syn_tsu113: string;
   attribute syn_tsu113 of DEF_ARCH : architecture is " F_FM0_ADDR[28]->CLK_BASE = 0.744";
   attribute syn_tsu114: string;
   attribute syn_tsu114 of DEF_ARCH : architecture is " F_FM0_ADDR[29]->CLK_BASE = 0.565";
   attribute syn_tsu115: string;
   attribute syn_tsu115 of DEF_ARCH : architecture is " F_FM0_ADDR[2]->CLK_BASE = 0.487";
   attribute syn_tsu116: string;
   attribute syn_tsu116 of DEF_ARCH : architecture is " F_FM0_ADDR[30]->CLK_BASE = 0.668";
   attribute syn_tsu117: string;
   attribute syn_tsu117 of DEF_ARCH : architecture is " F_FM0_ADDR[31]->CLK_BASE = 0.586";
   attribute syn_tsu118: string;
   attribute syn_tsu118 of DEF_ARCH : architecture is " F_FM0_ADDR[3]->CLK_BASE = 1.011";
   attribute syn_tsu119: string;
   attribute syn_tsu119 of DEF_ARCH : architecture is " F_FM0_ADDR[4]->CLK_BASE = 1.014";
   attribute syn_tsu120: string;
   attribute syn_tsu120 of DEF_ARCH : architecture is " F_FM0_ADDR[5]->CLK_BASE = 0.944";
   attribute syn_tsu121: string;
   attribute syn_tsu121 of DEF_ARCH : architecture is " F_FM0_ADDR[6]->CLK_BASE = 0.994";
   attribute syn_tsu122: string;
   attribute syn_tsu122 of DEF_ARCH : architecture is " F_FM0_ADDR[7]->CLK_BASE = 1.016";
   attribute syn_tsu123: string;
   attribute syn_tsu123 of DEF_ARCH : architecture is " F_FM0_ADDR[8]->CLK_BASE = 1.032";
   attribute syn_tsu124: string;
   attribute syn_tsu124 of DEF_ARCH : architecture is " F_FM0_ADDR[9]->CLK_BASE = 1.058";
   attribute syn_tsu125: string;
   attribute syn_tsu125 of DEF_ARCH : architecture is " F_FM0_ENABLE->CLK_BASE = 1.065";
   attribute syn_tsu126: string;
   attribute syn_tsu126 of DEF_ARCH : architecture is " F_FM0_SEL->CLK_BASE = 1.136";
   attribute syn_tsu127: string;
   attribute syn_tsu127 of DEF_ARCH : architecture is " F_FM0_WDATA[0]->CLK_BASE = 0.499";
   attribute syn_tsu128: string;
   attribute syn_tsu128 of DEF_ARCH : architecture is " F_FM0_WDATA[10]->CLK_BASE = 0.365";
   attribute syn_tsu129: string;
   attribute syn_tsu129 of DEF_ARCH : architecture is " F_FM0_WDATA[11]->CLK_BASE = 0.397";
   attribute syn_tsu130: string;
   attribute syn_tsu130 of DEF_ARCH : architecture is " F_FM0_WDATA[12]->CLK_BASE = 0.409";
   attribute syn_tsu131: string;
   attribute syn_tsu131 of DEF_ARCH : architecture is " F_FM0_WDATA[13]->CLK_BASE = 0.483";
   attribute syn_tsu132: string;
   attribute syn_tsu132 of DEF_ARCH : architecture is " F_FM0_WDATA[14]->CLK_BASE = 0.678";
   attribute syn_tsu133: string;
   attribute syn_tsu133 of DEF_ARCH : architecture is " F_FM0_WDATA[15]->CLK_BASE = 0.438";
   attribute syn_tsu134: string;
   attribute syn_tsu134 of DEF_ARCH : architecture is " F_FM0_WDATA[16]->CLK_BASE = 0.43";
   attribute syn_tsu135: string;
   attribute syn_tsu135 of DEF_ARCH : architecture is " F_FM0_WDATA[17]->CLK_BASE = 0.56";
   attribute syn_tsu136: string;
   attribute syn_tsu136 of DEF_ARCH : architecture is " F_FM0_WDATA[18]->CLK_BASE = 0.553";
   attribute syn_tsu137: string;
   attribute syn_tsu137 of DEF_ARCH : architecture is " F_FM0_WDATA[19]->CLK_BASE = 0.386";
   attribute syn_tsu138: string;
   attribute syn_tsu138 of DEF_ARCH : architecture is " F_FM0_WDATA[1]->CLK_BASE = 0.457";
   attribute syn_tsu139: string;
   attribute syn_tsu139 of DEF_ARCH : architecture is " F_FM0_WDATA[20]->CLK_BASE = 0.404";
   attribute syn_tsu140: string;
   attribute syn_tsu140 of DEF_ARCH : architecture is " F_FM0_WDATA[21]->CLK_BASE = 0.393";
   attribute syn_tsu141: string;
   attribute syn_tsu141 of DEF_ARCH : architecture is " F_FM0_WDATA[22]->CLK_BASE = 0.448";
   attribute syn_tsu142: string;
   attribute syn_tsu142 of DEF_ARCH : architecture is " F_FM0_WDATA[23]->CLK_BASE = 0.359";
   attribute syn_tsu143: string;
   attribute syn_tsu143 of DEF_ARCH : architecture is " F_FM0_WDATA[24]->CLK_BASE = 0.491";
   attribute syn_tsu144: string;
   attribute syn_tsu144 of DEF_ARCH : architecture is " F_FM0_WDATA[25]->CLK_BASE = 0.406";
   attribute syn_tsu145: string;
   attribute syn_tsu145 of DEF_ARCH : architecture is " F_FM0_WDATA[26]->CLK_BASE = 0.401";
   attribute syn_tsu146: string;
   attribute syn_tsu146 of DEF_ARCH : architecture is " F_FM0_WDATA[27]->CLK_BASE = 0.47";
   attribute syn_tsu147: string;
   attribute syn_tsu147 of DEF_ARCH : architecture is " F_FM0_WDATA[28]->CLK_BASE = 0.422";
   attribute syn_tsu148: string;
   attribute syn_tsu148 of DEF_ARCH : architecture is " F_FM0_WDATA[29]->CLK_BASE = 0.387";
   attribute syn_tsu149: string;
   attribute syn_tsu149 of DEF_ARCH : architecture is " F_FM0_WDATA[2]->CLK_BASE = 0.392";
   attribute syn_tsu150: string;
   attribute syn_tsu150 of DEF_ARCH : architecture is " F_FM0_WDATA[30]->CLK_BASE = 0.363";
   attribute syn_tsu151: string;
   attribute syn_tsu151 of DEF_ARCH : architecture is " F_FM0_WDATA[31]->CLK_BASE = 0.37";
   attribute syn_tsu152: string;
   attribute syn_tsu152 of DEF_ARCH : architecture is " F_FM0_WDATA[3]->CLK_BASE = 0.391";
   attribute syn_tsu153: string;
   attribute syn_tsu153 of DEF_ARCH : architecture is " F_FM0_WDATA[4]->CLK_BASE = 0.407";
   attribute syn_tsu154: string;
   attribute syn_tsu154 of DEF_ARCH : architecture is " F_FM0_WDATA[5]->CLK_BASE = 0.499";
   attribute syn_tsu155: string;
   attribute syn_tsu155 of DEF_ARCH : architecture is " F_FM0_WDATA[6]->CLK_BASE = 0.379";
   attribute syn_tsu156: string;
   attribute syn_tsu156 of DEF_ARCH : architecture is " F_FM0_WDATA[7]->CLK_BASE = 0.372";
   attribute syn_tsu157: string;
   attribute syn_tsu157 of DEF_ARCH : architecture is " F_FM0_WDATA[8]->CLK_BASE = 0.376";
   attribute syn_tsu158: string;
   attribute syn_tsu158 of DEF_ARCH : architecture is " F_FM0_WDATA[9]->CLK_BASE = 0.364";
   attribute syn_tsu159: string;
   attribute syn_tsu159 of DEF_ARCH : architecture is " F_FM0_WRITE->CLK_BASE = 0.569";
   attribute syn_tsu160: string;
   attribute syn_tsu160 of DEF_ARCH : architecture is " F_HM0_RDATA[0]->CLK_BASE = 0.357";
   attribute syn_tsu161: string;
   attribute syn_tsu161 of DEF_ARCH : architecture is " F_HM0_RDATA[10]->CLK_BASE = 0.37";
   attribute syn_tsu162: string;
   attribute syn_tsu162 of DEF_ARCH : architecture is " F_HM0_RDATA[11]->CLK_BASE = 0.393";
   attribute syn_tsu163: string;
   attribute syn_tsu163 of DEF_ARCH : architecture is " F_HM0_RDATA[12]->CLK_BASE = 0.522";
   attribute syn_tsu164: string;
   attribute syn_tsu164 of DEF_ARCH : architecture is " F_HM0_RDATA[13]->CLK_BASE = 0.312";
   attribute syn_tsu165: string;
   attribute syn_tsu165 of DEF_ARCH : architecture is " F_HM0_RDATA[14]->CLK_BASE = 0.344";
   attribute syn_tsu166: string;
   attribute syn_tsu166 of DEF_ARCH : architecture is " F_HM0_RDATA[15]->CLK_BASE = 0.355";
   attribute syn_tsu167: string;
   attribute syn_tsu167 of DEF_ARCH : architecture is " F_HM0_RDATA[16]->CLK_BASE = 0.409";
   attribute syn_tsu168: string;
   attribute syn_tsu168 of DEF_ARCH : architecture is " F_HM0_RDATA[17]->CLK_BASE = 0.467";
   attribute syn_tsu169: string;
   attribute syn_tsu169 of DEF_ARCH : architecture is " F_HM0_RDATA[18]->CLK_BASE = 0.466";
   attribute syn_tsu170: string;
   attribute syn_tsu170 of DEF_ARCH : architecture is " F_HM0_RDATA[19]->CLK_BASE = 0.31";
   attribute syn_tsu171: string;
   attribute syn_tsu171 of DEF_ARCH : architecture is " F_HM0_RDATA[1]->CLK_BASE = 0.445";
   attribute syn_tsu172: string;
   attribute syn_tsu172 of DEF_ARCH : architecture is " F_HM0_RDATA[20]->CLK_BASE = 0.333";
   attribute syn_tsu173: string;
   attribute syn_tsu173 of DEF_ARCH : architecture is " F_HM0_RDATA[21]->CLK_BASE = 0.404";
   attribute syn_tsu174: string;
   attribute syn_tsu174 of DEF_ARCH : architecture is " F_HM0_RDATA[22]->CLK_BASE = 0.423";
   attribute syn_tsu175: string;
   attribute syn_tsu175 of DEF_ARCH : architecture is " F_HM0_RDATA[23]->CLK_BASE = 0.432";
   attribute syn_tsu176: string;
   attribute syn_tsu176 of DEF_ARCH : architecture is " F_HM0_RDATA[24]->CLK_BASE = 0.342";
   attribute syn_tsu177: string;
   attribute syn_tsu177 of DEF_ARCH : architecture is " F_HM0_RDATA[25]->CLK_BASE = 0.386";
   attribute syn_tsu178: string;
   attribute syn_tsu178 of DEF_ARCH : architecture is " F_HM0_RDATA[26]->CLK_BASE = 0.335";
   attribute syn_tsu179: string;
   attribute syn_tsu179 of DEF_ARCH : architecture is " F_HM0_RDATA[27]->CLK_BASE = 0.374";
   attribute syn_tsu180: string;
   attribute syn_tsu180 of DEF_ARCH : architecture is " F_HM0_RDATA[28]->CLK_BASE = 0.434";
   attribute syn_tsu181: string;
   attribute syn_tsu181 of DEF_ARCH : architecture is " F_HM0_RDATA[29]->CLK_BASE = 0.43";
   attribute syn_tsu182: string;
   attribute syn_tsu182 of DEF_ARCH : architecture is " F_HM0_RDATA[2]->CLK_BASE = 0.34";
   attribute syn_tsu183: string;
   attribute syn_tsu183 of DEF_ARCH : architecture is " F_HM0_RDATA[30]->CLK_BASE = 0.419";
   attribute syn_tsu184: string;
   attribute syn_tsu184 of DEF_ARCH : architecture is " F_HM0_RDATA[31]->CLK_BASE = 0.441";
   attribute syn_tsu185: string;
   attribute syn_tsu185 of DEF_ARCH : architecture is " F_HM0_RDATA[3]->CLK_BASE = 0.351";
   attribute syn_tsu186: string;
   attribute syn_tsu186 of DEF_ARCH : architecture is " F_HM0_RDATA[4]->CLK_BASE = 0.376";
   attribute syn_tsu187: string;
   attribute syn_tsu187 of DEF_ARCH : architecture is " F_HM0_RDATA[5]->CLK_BASE = 0.433";
   attribute syn_tsu188: string;
   attribute syn_tsu188 of DEF_ARCH : architecture is " F_HM0_RDATA[6]->CLK_BASE = 0.379";
   attribute syn_tsu189: string;
   attribute syn_tsu189 of DEF_ARCH : architecture is " F_HM0_RDATA[7]->CLK_BASE = 0.357";
   attribute syn_tsu190: string;
   attribute syn_tsu190 of DEF_ARCH : architecture is " F_HM0_RDATA[8]->CLK_BASE = 0.374";
   attribute syn_tsu191: string;
   attribute syn_tsu191 of DEF_ARCH : architecture is " F_HM0_RDATA[9]->CLK_BASE = 0.352";
   attribute syn_tsu192: string;
   attribute syn_tsu192 of DEF_ARCH : architecture is " F_HM0_READY->CLK_BASE = 1.559";
   attribute syn_tsu193: string;
   attribute syn_tsu193 of DEF_ARCH : architecture is " F_HM0_RESP->CLK_BASE = 0.895";
   attribute syn_tsu194: string;
   attribute syn_tsu194 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[0]->CLK_BASE = 1.188";
   attribute syn_tsu195: string;
   attribute syn_tsu195 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[10]->CLK_BASE = 0.452";
   attribute syn_tsu196: string;
   attribute syn_tsu196 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[11]->CLK_BASE = 0.688";
   attribute syn_tsu197: string;
   attribute syn_tsu197 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[12]->CLK_BASE = 0.601";
   attribute syn_tsu198: string;
   attribute syn_tsu198 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[13]->CLK_BASE = 0.605";
   attribute syn_tsu199: string;
   attribute syn_tsu199 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[14]->CLK_BASE = 0.576";
   attribute syn_tsu200: string;
   attribute syn_tsu200 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[15]->CLK_BASE = 0.662";
   attribute syn_tsu201: string;
   attribute syn_tsu201 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[16]->CLK_BASE = 0.421";
   attribute syn_tsu202: string;
   attribute syn_tsu202 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[17]->CLK_BASE = 0.584";
   attribute syn_tsu203: string;
   attribute syn_tsu203 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[18]->CLK_BASE = 0.65";
   attribute syn_tsu204: string;
   attribute syn_tsu204 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[19]->CLK_BASE = 0.928";
   attribute syn_tsu205: string;
   attribute syn_tsu205 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[1]->CLK_BASE = 1.161";
   attribute syn_tsu206: string;
   attribute syn_tsu206 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[20]->CLK_BASE = 0.743";
   attribute syn_tsu207: string;
   attribute syn_tsu207 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[21]->CLK_BASE = 0.643";
   attribute syn_tsu208: string;
   attribute syn_tsu208 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[22]->CLK_BASE = 0.597";
   attribute syn_tsu209: string;
   attribute syn_tsu209 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[23]->CLK_BASE = 0.537";
   attribute syn_tsu210: string;
   attribute syn_tsu210 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[24]->CLK_BASE = 0.695";
   attribute syn_tsu211: string;
   attribute syn_tsu211 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[25]->CLK_BASE = 0.592";
   attribute syn_tsu212: string;
   attribute syn_tsu212 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[26]->CLK_BASE = 0.552";
   attribute syn_tsu213: string;
   attribute syn_tsu213 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[27]->CLK_BASE = 0.591";
   attribute syn_tsu214: string;
   attribute syn_tsu214 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[28]->CLK_BASE = 0.586";
   attribute syn_tsu215: string;
   attribute syn_tsu215 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[29]->CLK_BASE = 0.563";
   attribute syn_tsu216: string;
   attribute syn_tsu216 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[2]->CLK_BASE = 1.281";
   attribute syn_tsu217: string;
   attribute syn_tsu217 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[30]->CLK_BASE = 0.437";
   attribute syn_tsu218: string;
   attribute syn_tsu218 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[31]->CLK_BASE = 0.633";
   attribute syn_tsu219: string;
   attribute syn_tsu219 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[32]->CLK_BASE = 0.805";
   attribute syn_tsu220: string;
   attribute syn_tsu220 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[33]->CLK_BASE = 0.992";
   attribute syn_tsu221: string;
   attribute syn_tsu221 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[34]->CLK_BASE = 0.945";
   attribute syn_tsu222: string;
   attribute syn_tsu222 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[35]->CLK_BASE = 1.244";
   attribute syn_tsu223: string;
   attribute syn_tsu223 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[36]->CLK_BASE = 0.82";
   attribute syn_tsu224: string;
   attribute syn_tsu224 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[37]->CLK_BASE = 1.218";
   attribute syn_tsu225: string;
   attribute syn_tsu225 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[38]->CLK_BASE = 1.179";
   attribute syn_tsu226: string;
   attribute syn_tsu226 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[39]->CLK_BASE = 0.945";
   attribute syn_tsu227: string;
   attribute syn_tsu227 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[3]->CLK_BASE = 1.301";
   attribute syn_tsu228: string;
   attribute syn_tsu228 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[40]->CLK_BASE = 0.732";
   attribute syn_tsu229: string;
   attribute syn_tsu229 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[41]->CLK_BASE = 0.602";
   attribute syn_tsu230: string;
   attribute syn_tsu230 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[42]->CLK_BASE = 0.5";
   attribute syn_tsu231: string;
   attribute syn_tsu231 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[43]->CLK_BASE = 0.647";
   attribute syn_tsu232: string;
   attribute syn_tsu232 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[44]->CLK_BASE = 0.695";
   attribute syn_tsu233: string;
   attribute syn_tsu233 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[45]->CLK_BASE = 0.766";
   attribute syn_tsu234: string;
   attribute syn_tsu234 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[46]->CLK_BASE = 0.641";
   attribute syn_tsu235: string;
   attribute syn_tsu235 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[47]->CLK_BASE = 0.66";
   attribute syn_tsu236: string;
   attribute syn_tsu236 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[48]->CLK_BASE = 0.587";
   attribute syn_tsu237: string;
   attribute syn_tsu237 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[49]->CLK_BASE = 0.738";
   attribute syn_tsu238: string;
   attribute syn_tsu238 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[4]->CLK_BASE = 0.946";
   attribute syn_tsu239: string;
   attribute syn_tsu239 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[50]->CLK_BASE = 0.614";
   attribute syn_tsu240: string;
   attribute syn_tsu240 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[51]->CLK_BASE = 0.72";
   attribute syn_tsu241: string;
   attribute syn_tsu241 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[52]->CLK_BASE = 0.482";
   attribute syn_tsu242: string;
   attribute syn_tsu242 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[53]->CLK_BASE = 0.782";
   attribute syn_tsu243: string;
   attribute syn_tsu243 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[54]->CLK_BASE = 0.635";
   attribute syn_tsu244: string;
   attribute syn_tsu244 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[55]->CLK_BASE = 0.579";
   attribute syn_tsu245: string;
   attribute syn_tsu245 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[56]->CLK_BASE = 0.604";
   attribute syn_tsu246: string;
   attribute syn_tsu246 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[57]->CLK_BASE = 0.704";
   attribute syn_tsu247: string;
   attribute syn_tsu247 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[58]->CLK_BASE = 0.459";
   attribute syn_tsu248: string;
   attribute syn_tsu248 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[59]->CLK_BASE = 0.888";
   attribute syn_tsu249: string;
   attribute syn_tsu249 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[5]->CLK_BASE = 0.863";
   attribute syn_tsu250: string;
   attribute syn_tsu250 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[60]->CLK_BASE = 0.554";
   attribute syn_tsu251: string;
   attribute syn_tsu251 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[61]->CLK_BASE = 0.517";
   attribute syn_tsu252: string;
   attribute syn_tsu252 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[62]->CLK_BASE = 0.69";
   attribute syn_tsu253: string;
   attribute syn_tsu253 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[63]->CLK_BASE = 0.618";
   attribute syn_tsu254: string;
   attribute syn_tsu254 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[6]->CLK_BASE = 1.142";
   attribute syn_tsu255: string;
   attribute syn_tsu255 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[7]->CLK_BASE = 1.188";
   attribute syn_tsu256: string;
   attribute syn_tsu256 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[8]->CLK_BASE = 0.61";
   attribute syn_tsu257: string;
   attribute syn_tsu257 of DEF_ARCH : architecture is " F_WDATA_HWDATA01[9]->CLK_BASE = 0.774";
   attribute syn_tsu258: string;
   attribute syn_tsu258 of DEF_ARCH : architecture is " F_WID_HREADY01[0]->CLK_BASE = 1.93";
   attribute syn_tsu259: string;
   attribute syn_tsu259 of DEF_ARCH : architecture is " F_WID_HREADY01[1]->CLK_BASE = 1.571";
   attribute syn_tsu260: string;
   attribute syn_tsu260 of DEF_ARCH : architecture is " F_WLAST->CLK_BASE = 1.039";
   attribute syn_tsu261: string;
   attribute syn_tsu261 of DEF_ARCH : architecture is " I2C0_SDA_F2H_SCP->I2C0_SCL_F2H_SCP = 0.197";
   attribute syn_tsu262: string;
   attribute syn_tsu262 of DEF_ARCH : architecture is " I2C1_SDA_F2H_SCP->I2C1_SCL_F2H_SCP = 0.279";
   attribute syn_tsu263: string;
   attribute syn_tsu263 of DEF_ARCH : architecture is " MGPIO0A_F2H_GPIN->CLK_BASE = 0.626";
   attribute syn_tsu264: string;
   attribute syn_tsu264 of DEF_ARCH : architecture is " MGPIO11B_F2H_GPIN->CLK_BASE = 0.603";
   attribute syn_tsu265: string;
   attribute syn_tsu265 of DEF_ARCH : architecture is " MGPIO17B_F2H_GPIN->CLK_BASE = 0.561";
   attribute syn_tsu266: string;
   attribute syn_tsu266 of DEF_ARCH : architecture is " MGPIO18B_F2H_GPIN->CLK_BASE = 0.694";
   attribute syn_tsu267: string;
   attribute syn_tsu267 of DEF_ARCH : architecture is " MGPIO24B_F2H_GPIN->CLK_BASE = 0.568";
   attribute syn_tsu268: string;
   attribute syn_tsu268 of DEF_ARCH : architecture is " MGPIO27B_F2H_GPIN->CLK_BASE = 0.655";
   attribute syn_tsu269: string;
   attribute syn_tsu269 of DEF_ARCH : architecture is " MGPIO28B_F2H_GPIN->CLK_BASE = 0.732";
   attribute syn_tsu270: string;
   attribute syn_tsu270 of DEF_ARCH : architecture is " MGPIO2A_F2H_GPIN->CLK_BASE = 0.666";
   attribute syn_tsu271: string;
   attribute syn_tsu271 of DEF_ARCH : architecture is " MGPIO30B_F2H_GPIN->CLK_BASE = 0.659";
   attribute syn_tsu272: string;
   attribute syn_tsu272 of DEF_ARCH : architecture is " MGPIO31B_F2H_GPIN->CLK_BASE = 0.83";
   attribute syn_tsu273: string;
   attribute syn_tsu273 of DEF_ARCH : architecture is " MGPIO3A_F2H_GPIN->CLK_BASE = 0.547";
   attribute syn_tsu274: string;
   attribute syn_tsu274 of DEF_ARCH : architecture is " MGPIO4A_F2H_GPIN->CLK_BASE = 0.784";
   attribute syn_tsu275: string;
   attribute syn_tsu275 of DEF_ARCH : architecture is " MGPIO5A_F2H_GPIN->CLK_BASE = 0.706";
   attribute syn_tsu276: string;
   attribute syn_tsu276 of DEF_ARCH : architecture is " MGPIO6A_F2H_GPIN->CLK_BASE = 0.593";
   attribute syn_tsu277: string;
   attribute syn_tsu277 of DEF_ARCH : architecture is " MGPIO7A_F2H_GPIN->CLK_BASE = 0.64";
   attribute syn_tsu278: string;
   attribute syn_tsu278 of DEF_ARCH : architecture is " MMUART0_CTS_F2H_SCP->CLK_BASE = 1.146";
   attribute syn_tsu279: string;
   attribute syn_tsu279 of DEF_ARCH : architecture is " MMUART0_DCD_F2H_SCP->CLK_BASE = 1.219";
   attribute syn_tsu280: string;
   attribute syn_tsu280 of DEF_ARCH : architecture is " MMUART0_DSR_F2H_SCP->CLK_BASE = 1.17";
   attribute syn_tsu281: string;
   attribute syn_tsu281 of DEF_ARCH : architecture is " MMUART0_RI_F2H_SCP->CLK_BASE = 0.83";
   attribute syn_tsu282: string;
   attribute syn_tsu282 of DEF_ARCH : architecture is " MMUART0_SCK_F2H_SCP->CLK_BASE = 1.081";
   attribute syn_tsu283: string;
   attribute syn_tsu283 of DEF_ARCH : architecture is " MMUART0_TXD_F2H_SCP->CLK_BASE = 1.216";
   attribute syn_tsu284: string;
   attribute syn_tsu284 of DEF_ARCH : architecture is " MMUART1_CTS_F2H_SCP->CLK_BASE = 1.062";
   attribute syn_tsu285: string;
   attribute syn_tsu285 of DEF_ARCH : architecture is " MMUART1_DCD_F2H_SCP->CLK_BASE = 0.933";
   attribute syn_tsu286: string;
   attribute syn_tsu286 of DEF_ARCH : architecture is " MMUART1_DSR_F2H_SCP->CLK_BASE = 1.021";
   attribute syn_tsu287: string;
   attribute syn_tsu287 of DEF_ARCH : architecture is " MMUART1_RI_F2H_SCP->CLK_BASE = 0.822";
   attribute syn_tsu288: string;
   attribute syn_tsu288 of DEF_ARCH : architecture is " MMUART1_RXD_F2H_SCP->CLK_BASE = 1.186";
   attribute syn_tsu289: string;
   attribute syn_tsu289 of DEF_ARCH : architecture is " MMUART1_SCK_F2H_SCP->CLK_BASE = 0.811";
   attribute syn_tsu290: string;
   attribute syn_tsu290 of DEF_ARCH : architecture is " MMUART1_TXD_F2H_SCP->CLK_BASE = 1.064";
   attribute syn_tsu291: string;
   attribute syn_tsu291 of DEF_ARCH : architecture is " SMBALERT_NI0->I2C0_SCL_F2H_SCP = 0";
   attribute syn_tsu292: string;
   attribute syn_tsu292 of DEF_ARCH : architecture is " SMBALERT_NI1->I2C1_SCL_F2H_SCP = 0";
   attribute syn_tsu293: string;
   attribute syn_tsu293 of DEF_ARCH : architecture is " SMBSUS_NI0->I2C0_SCL_F2H_SCP = 0";
   attribute syn_tsu294: string;
   attribute syn_tsu294 of DEF_ARCH : architecture is " SMBSUS_NI1->I2C1_SCL_F2H_SCP = 0";
   attribute syn_tsu295: string;
   attribute syn_tsu295 of DEF_ARCH : architecture is " SPI1_SDI_F2H_SCP->SPI1_CLK_IN = 1.206";
   attribute syn_tco0: string;
   attribute syn_tco0 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_A = 3.439";
   attribute syn_tco1: string;
   attribute syn_tco1 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_B = 3.465";
   attribute syn_tco2: string;
   attribute syn_tco2 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_A = 3.364";
   attribute syn_tco3: string;
   attribute syn_tco3 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_B = 3.451";
   attribute syn_tco4: string;
   attribute syn_tco4 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT = 3.846";
   attribute syn_tco5: string;
   attribute syn_tco5 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_A = 3.438";
   attribute syn_tco6: string;
   attribute syn_tco6 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_B = 3.340";
   attribute syn_tco7: string;
   attribute syn_tco7 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT = 3.752";
   attribute syn_tco8: string;
   attribute syn_tco8 of DEF_ARCH : architecture is " CLK_BASE->F_ARREADY_HREADYOUT1 = 3.673";
   attribute syn_tco9: string;
   attribute syn_tco9 of DEF_ARCH : architecture is " CLK_BASE->F_BID[0] = 3.895";
   attribute syn_tco10: string;
   attribute syn_tco10 of DEF_ARCH : architecture is " CLK_BASE->F_BID[1] = 3.893";
   attribute syn_tco11: string;
   attribute syn_tco11 of DEF_ARCH : architecture is " CLK_BASE->F_BID[2] = 3.968";
   attribute syn_tco12: string;
   attribute syn_tco12 of DEF_ARCH : architecture is " CLK_BASE->F_BRESP_HRESP0[0] = 4.343";
   attribute syn_tco13: string;
   attribute syn_tco13 of DEF_ARCH : architecture is " CLK_BASE->F_BRESP_HRESP0[1] = 4.945";
   attribute syn_tco14: string;
   attribute syn_tco14 of DEF_ARCH : architecture is " CLK_BASE->F_BVALID = 3.969";
   attribute syn_tco15: string;
   attribute syn_tco15 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[0] = 4.297";
   attribute syn_tco16: string;
   attribute syn_tco16 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[10] = 4.255";
   attribute syn_tco17: string;
   attribute syn_tco17 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[11] = 4.154";
   attribute syn_tco18: string;
   attribute syn_tco18 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[12] = 4.326";
   attribute syn_tco19: string;
   attribute syn_tco19 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[13] = 4.327";
   attribute syn_tco20: string;
   attribute syn_tco20 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[14] = 4.205";
   attribute syn_tco21: string;
   attribute syn_tco21 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[15] = 4.159";
   attribute syn_tco22: string;
   attribute syn_tco22 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[16] = 4.240";
   attribute syn_tco23: string;
   attribute syn_tco23 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[17] = 4.244";
   attribute syn_tco24: string;
   attribute syn_tco24 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[18] = 4.216";
   attribute syn_tco25: string;
   attribute syn_tco25 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[19] = 4.246";
   attribute syn_tco26: string;
   attribute syn_tco26 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[1] = 4.187";
   attribute syn_tco27: string;
   attribute syn_tco27 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[20] = 4.281";
   attribute syn_tco28: string;
   attribute syn_tco28 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[21] = 4.277";
   attribute syn_tco29: string;
   attribute syn_tco29 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[22] = 4.240";
   attribute syn_tco30: string;
   attribute syn_tco30 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[23] = 4.230";
   attribute syn_tco31: string;
   attribute syn_tco31 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[24] = 4.272";
   attribute syn_tco32: string;
   attribute syn_tco32 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[25] = 4.259";
   attribute syn_tco33: string;
   attribute syn_tco33 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[26] = 4.225";
   attribute syn_tco34: string;
   attribute syn_tco34 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[27] = 4.316";
   attribute syn_tco35: string;
   attribute syn_tco35 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[28] = 4.274";
   attribute syn_tco36: string;
   attribute syn_tco36 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[29] = 4.293";
   attribute syn_tco37: string;
   attribute syn_tco37 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[2] = 4.281";
   attribute syn_tco38: string;
   attribute syn_tco38 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[30] = 4.190";
   attribute syn_tco39: string;
   attribute syn_tco39 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[31] = 4.206";
   attribute syn_tco40: string;
   attribute syn_tco40 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[3] = 4.304";
   attribute syn_tco41: string;
   attribute syn_tco41 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[4] = 4.240";
   attribute syn_tco42: string;
   attribute syn_tco42 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[5] = 4.160";
   attribute syn_tco43: string;
   attribute syn_tco43 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[6] = 4.123";
   attribute syn_tco44: string;
   attribute syn_tco44 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[7] = 4.168";
   attribute syn_tco45: string;
   attribute syn_tco45 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[8] = 4.245";
   attribute syn_tco46: string;
   attribute syn_tco46 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[9] = 4.141";
   attribute syn_tco47: string;
   attribute syn_tco47 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_READYOUT = 3.950";
   attribute syn_tco48: string;
   attribute syn_tco48 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RESP = 3.881";
   attribute syn_tco49: string;
   attribute syn_tco49 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[0] = 3.467";
   attribute syn_tco50: string;
   attribute syn_tco50 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[10] = 3.247";
   attribute syn_tco51: string;
   attribute syn_tco51 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[11] = 3.262";
   attribute syn_tco52: string;
   attribute syn_tco52 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[12] = 3.203";
   attribute syn_tco53: string;
   attribute syn_tco53 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[13] = 3.243";
   attribute syn_tco54: string;
   attribute syn_tco54 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[14] = 3.210";
   attribute syn_tco55: string;
   attribute syn_tco55 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[15] = 3.237";
   attribute syn_tco56: string;
   attribute syn_tco56 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[16] = 3.254";
   attribute syn_tco57: string;
   attribute syn_tco57 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[17] = 3.250";
   attribute syn_tco58: string;
   attribute syn_tco58 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[18] = 3.238";
   attribute syn_tco59: string;
   attribute syn_tco59 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[19] = 3.226";
   attribute syn_tco60: string;
   attribute syn_tco60 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[1] = 3.508";
   attribute syn_tco61: string;
   attribute syn_tco61 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[20] = 3.219";
   attribute syn_tco62: string;
   attribute syn_tco62 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[21] = 3.222";
   attribute syn_tco63: string;
   attribute syn_tco63 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[22] = 3.244";
   attribute syn_tco64: string;
   attribute syn_tco64 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[23] = 3.277";
   attribute syn_tco65: string;
   attribute syn_tco65 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[24] = 3.194";
   attribute syn_tco66: string;
   attribute syn_tco66 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[25] = 3.228";
   attribute syn_tco67: string;
   attribute syn_tco67 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[26] = 3.270";
   attribute syn_tco68: string;
   attribute syn_tco68 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[27] = 3.226";
   attribute syn_tco69: string;
   attribute syn_tco69 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[28] = 3.261";
   attribute syn_tco70: string;
   attribute syn_tco70 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[29] = 3.191";
   attribute syn_tco71: string;
   attribute syn_tco71 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[2] = 3.266";
   attribute syn_tco72: string;
   attribute syn_tco72 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[30] = 3.225";
   attribute syn_tco73: string;
   attribute syn_tco73 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[31] = 3.261";
   attribute syn_tco74: string;
   attribute syn_tco74 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[3] = 3.231";
   attribute syn_tco75: string;
   attribute syn_tco75 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[4] = 3.236";
   attribute syn_tco76: string;
   attribute syn_tco76 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[5] = 3.253";
   attribute syn_tco77: string;
   attribute syn_tco77 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[6] = 3.234";
   attribute syn_tco78: string;
   attribute syn_tco78 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[7] = 3.222";
   attribute syn_tco79: string;
   attribute syn_tco79 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[8] = 3.275";
   attribute syn_tco80: string;
   attribute syn_tco80 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[9] = 3.222";
   attribute syn_tco81: string;
   attribute syn_tco81 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ENABLE = 3.399";
   attribute syn_tco82: string;
   attribute syn_tco82 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SEL = 3.297";
   attribute syn_tco83: string;
   attribute syn_tco83 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[0] = 3.200";
   attribute syn_tco84: string;
   attribute syn_tco84 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[10] = 3.343";
   attribute syn_tco85: string;
   attribute syn_tco85 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[11] = 3.396";
   attribute syn_tco86: string;
   attribute syn_tco86 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[12] = 3.330";
   attribute syn_tco87: string;
   attribute syn_tco87 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[13] = 3.479";
   attribute syn_tco88: string;
   attribute syn_tco88 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[14] = 3.261";
   attribute syn_tco89: string;
   attribute syn_tco89 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[15] = 3.391";
   attribute syn_tco90: string;
   attribute syn_tco90 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[16] = 3.362";
   attribute syn_tco91: string;
   attribute syn_tco91 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[17] = 3.406";
   attribute syn_tco92: string;
   attribute syn_tco92 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[18] = 3.333";
   attribute syn_tco93: string;
   attribute syn_tco93 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[19] = 3.466";
   attribute syn_tco94: string;
   attribute syn_tco94 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[1] = 3.207";
   attribute syn_tco95: string;
   attribute syn_tco95 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[20] = 3.335";
   attribute syn_tco96: string;
   attribute syn_tco96 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[21] = 3.457";
   attribute syn_tco97: string;
   attribute syn_tco97 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[22] = 3.420";
   attribute syn_tco98: string;
   attribute syn_tco98 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[23] = 3.129";
   attribute syn_tco99: string;
   attribute syn_tco99 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[24] = 3.325";
   attribute syn_tco100: string;
   attribute syn_tco100 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[25] = 3.482";
   attribute syn_tco101: string;
   attribute syn_tco101 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[26] = 3.516";
   attribute syn_tco102: string;
   attribute syn_tco102 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[27] = 3.480";
   attribute syn_tco103: string;
   attribute syn_tco103 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[28] = 3.453";
   attribute syn_tco104: string;
   attribute syn_tco104 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[29] = 3.514";
   attribute syn_tco105: string;
   attribute syn_tco105 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[2] = 3.287";
   attribute syn_tco106: string;
   attribute syn_tco106 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[30] = 3.565";
   attribute syn_tco107: string;
   attribute syn_tco107 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[31] = 3.516";
   attribute syn_tco108: string;
   attribute syn_tco108 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[3] = 3.144";
   attribute syn_tco109: string;
   attribute syn_tco109 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[4] = 3.342";
   attribute syn_tco110: string;
   attribute syn_tco110 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[5] = 3.331";
   attribute syn_tco111: string;
   attribute syn_tco111 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[6] = 3.421";
   attribute syn_tco112: string;
   attribute syn_tco112 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[7] = 3.428";
   attribute syn_tco113: string;
   attribute syn_tco113 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[8] = 3.434";
   attribute syn_tco114: string;
   attribute syn_tco114 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[9] = 3.423";
   attribute syn_tco115: string;
   attribute syn_tco115 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WRITE = 3.634";
   attribute syn_tco116: string;
   attribute syn_tco116 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[0] = 3.872";
   attribute syn_tco117: string;
   attribute syn_tco117 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[10] = 3.924";
   attribute syn_tco118: string;
   attribute syn_tco118 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[11] = 4.030";
   attribute syn_tco119: string;
   attribute syn_tco119 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[12] = 4.007";
   attribute syn_tco120: string;
   attribute syn_tco120 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[13] = 4.058";
   attribute syn_tco121: string;
   attribute syn_tco121 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[14] = 4.246";
   attribute syn_tco122: string;
   attribute syn_tco122 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[15] = 4.084";
   attribute syn_tco123: string;
   attribute syn_tco123 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[16] = 4.202";
   attribute syn_tco124: string;
   attribute syn_tco124 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[17] = 4.073";
   attribute syn_tco125: string;
   attribute syn_tco125 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[18] = 4.169";
   attribute syn_tco126: string;
   attribute syn_tco126 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[19] = 3.988";
   attribute syn_tco127: string;
   attribute syn_tco127 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[1] = 3.877";
   attribute syn_tco128: string;
   attribute syn_tco128 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[20] = 4.099";
   attribute syn_tco129: string;
   attribute syn_tco129 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[21] = 3.921";
   attribute syn_tco130: string;
   attribute syn_tco130 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[22] = 3.693";
   attribute syn_tco131: string;
   attribute syn_tco131 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[23] = 4.061";
   attribute syn_tco132: string;
   attribute syn_tco132 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[24] = 3.879";
   attribute syn_tco133: string;
   attribute syn_tco133 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[25] = 3.960";
   attribute syn_tco134: string;
   attribute syn_tco134 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[26] = 4.019";
   attribute syn_tco135: string;
   attribute syn_tco135 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[27] = 3.932";
   attribute syn_tco136: string;
   attribute syn_tco136 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[28] = 4.105";
   attribute syn_tco137: string;
   attribute syn_tco137 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[29] = 3.830";
   attribute syn_tco138: string;
   attribute syn_tco138 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[2] = 4.115";
   attribute syn_tco139: string;
   attribute syn_tco139 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[30] = 3.857";
   attribute syn_tco140: string;
   attribute syn_tco140 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[31] = 3.837";
   attribute syn_tco141: string;
   attribute syn_tco141 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[32] = 4.083";
   attribute syn_tco142: string;
   attribute syn_tco142 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[33] = 3.910";
   attribute syn_tco143: string;
   attribute syn_tco143 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[34] = 3.967";
   attribute syn_tco144: string;
   attribute syn_tco144 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[35] = 3.929";
   attribute syn_tco145: string;
   attribute syn_tco145 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[36] = 3.983";
   attribute syn_tco146: string;
   attribute syn_tco146 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[37] = 4.158";
   attribute syn_tco147: string;
   attribute syn_tco147 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[38] = 4.327";
   attribute syn_tco148: string;
   attribute syn_tco148 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[39] = 4.221";
   attribute syn_tco149: string;
   attribute syn_tco149 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[3] = 4.100";
   attribute syn_tco150: string;
   attribute syn_tco150 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[40] = 3.917";
   attribute syn_tco151: string;
   attribute syn_tco151 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[41] = 3.937";
   attribute syn_tco152: string;
   attribute syn_tco152 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[42] = 3.911";
   attribute syn_tco153: string;
   attribute syn_tco153 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[43] = 3.782";
   attribute syn_tco154: string;
   attribute syn_tco154 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[44] = 4.063";
   attribute syn_tco155: string;
   attribute syn_tco155 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[45] = 4.203";
   attribute syn_tco156: string;
   attribute syn_tco156 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[46] = 3.913";
   attribute syn_tco157: string;
   attribute syn_tco157 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[47] = 3.970";
   attribute syn_tco158: string;
   attribute syn_tco158 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[48] = 3.715";
   attribute syn_tco159: string;
   attribute syn_tco159 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[49] = 3.845";
   attribute syn_tco160: string;
   attribute syn_tco160 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[4] = 4.013";
   attribute syn_tco161: string;
   attribute syn_tco161 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[50] = 4.033";
   attribute syn_tco162: string;
   attribute syn_tco162 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[51] = 4.282";
   attribute syn_tco163: string;
   attribute syn_tco163 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[52] = 4.329";
   attribute syn_tco164: string;
   attribute syn_tco164 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[53] = 3.969";
   attribute syn_tco165: string;
   attribute syn_tco165 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[54] = 3.908";
   attribute syn_tco166: string;
   attribute syn_tco166 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[55] = 3.927";
   attribute syn_tco167: string;
   attribute syn_tco167 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[56] = 4.309";
   attribute syn_tco168: string;
   attribute syn_tco168 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[57] = 4.360";
   attribute syn_tco169: string;
   attribute syn_tco169 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[58] = 4.123";
   attribute syn_tco170: string;
   attribute syn_tco170 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[59] = 4.086";
   attribute syn_tco171: string;
   attribute syn_tco171 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[5] = 4.131";
   attribute syn_tco172: string;
   attribute syn_tco172 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[60] = 4.055";
   attribute syn_tco173: string;
   attribute syn_tco173 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[61] = 4.245";
   attribute syn_tco174: string;
   attribute syn_tco174 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[62] = 4.075";
   attribute syn_tco175: string;
   attribute syn_tco175 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[63] = 3.868";
   attribute syn_tco176: string;
   attribute syn_tco176 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[6] = 4.052";
   attribute syn_tco177: string;
   attribute syn_tco177 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[7] = 3.936";
   attribute syn_tco178: string;
   attribute syn_tco178 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[8] = 3.883";
   attribute syn_tco179: string;
   attribute syn_tco179 of DEF_ARCH : architecture is " CLK_BASE->F_RDATA_HRDATA01[9] = 4.177";
   attribute syn_tco180: string;
   attribute syn_tco180 of DEF_ARCH : architecture is " CLK_BASE->F_RID[0] = 4.070";
   attribute syn_tco181: string;
   attribute syn_tco181 of DEF_ARCH : architecture is " CLK_BASE->F_RID[1] = 3.915";
   attribute syn_tco182: string;
   attribute syn_tco182 of DEF_ARCH : architecture is " CLK_BASE->F_RRESP_HRESP1[0] = 3.775";
   attribute syn_tco183: string;
   attribute syn_tco183 of DEF_ARCH : architecture is " CLK_BASE->H2FCALIB = 3.131";
   attribute syn_tco184: string;
   attribute syn_tco184 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_MGPIO31B_H2F_B = 3.495";
   attribute syn_tco185: string;
   attribute syn_tco185 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_USBC_DATA1_MGPIO31B_OE = 3.495";
   attribute syn_tco186: string;
   attribute syn_tco186 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_A = 3.541";
   attribute syn_tco187: string;
   attribute syn_tco187 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_B = 3.437";
   attribute syn_tco188: string;
   attribute syn_tco188 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_USBC_DATA0_MGPIO30B_OE = 2.923";
   attribute syn_tco189: string;
   attribute syn_tco189 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_MGPIO1A_H2F_B = 3.445";
   attribute syn_tco190: string;
   attribute syn_tco190 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OE = 2.802";
   attribute syn_tco191: string;
   attribute syn_tco191 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OUT = 3.792";
   attribute syn_tco192: string;
   attribute syn_tco192 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_A = 3.387";
   attribute syn_tco193: string;
   attribute syn_tco193 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_B = 3.538";
   attribute syn_tco194: string;
   attribute syn_tco194 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_USBA_DATA3_MGPIO0A_OE = 3.370";
   attribute syn_tco195: string;
   attribute syn_tco195 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OE = 2.823";
   attribute syn_tco196: string;
   attribute syn_tco196 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OUT = 2.743";
   attribute syn_tco197: string;
   attribute syn_tco197 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OE = 2.781";
   attribute syn_tco198: string;
   attribute syn_tco198 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OUT = 2.864";
   attribute syn_tco199: string;
   attribute syn_tco199 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_A = 3.403";
   attribute syn_tco200: string;
   attribute syn_tco200 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_B = 3.548";
   attribute syn_tco201: string;
   attribute syn_tco201 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_USBC_DATA7_MGPIO19B_OE = 3.197";
   attribute syn_tco202: string;
   attribute syn_tco202 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT = 3.548";
   attribute syn_tco203: string;
   attribute syn_tco203 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_A = 3.267";
   attribute syn_tco204: string;
   attribute syn_tco204 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_B = 3.437";
   attribute syn_tco205: string;
   attribute syn_tco205 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_OE = 2.977";
   attribute syn_tco206: string;
   attribute syn_tco206 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_OUT = 3.318";
   attribute syn_tco207: string;
   attribute syn_tco207 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_A = 3.295";
   attribute syn_tco208: string;
   attribute syn_tco208 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_B = 3.486";
   attribute syn_tco209: string;
   attribute syn_tco209 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_OE = 2.994";
   attribute syn_tco210: string;
   attribute syn_tco210 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_OUT = 3.371";
   attribute syn_tco211: string;
   attribute syn_tco211 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_A = 3.273";
   attribute syn_tco212: string;
   attribute syn_tco212 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_B = 3.403";
   attribute syn_tco213: string;
   attribute syn_tco213 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT = 2.864";
   attribute syn_tco214: string;
   attribute syn_tco214 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_A = 3.493";
   attribute syn_tco215: string;
   attribute syn_tco215 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_B = 3.454";
   attribute syn_tco216: string;
   attribute syn_tco216 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_OE = 3.278";
   attribute syn_tco217: string;
   attribute syn_tco217 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_OUT = 2.887";
   attribute syn_tco218: string;
   attribute syn_tco218 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_A = 3.483";
   attribute syn_tco219: string;
   attribute syn_tco219 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_B = 3.441";
   attribute syn_tco220: string;
   attribute syn_tco220 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT = 2.981";
   attribute syn_tco221: string;
   attribute syn_tco221 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_A = 3.548";
   attribute syn_tco222: string;
   attribute syn_tco222 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_B = 3.469";
   attribute syn_tco223: string;
   attribute syn_tco223 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_A = 3.323";
   attribute syn_tco224: string;
   attribute syn_tco224 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_B = 3.442";
   attribute syn_tco225: string;
   attribute syn_tco225 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OE = 3.085";
   attribute syn_tco226: string;
   attribute syn_tco226 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OUT = 3.061";
   attribute syn_tco227: string;
   attribute syn_tco227 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_A = 3.541";
   attribute syn_tco228: string;
   attribute syn_tco228 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_B = 3.439";
   attribute syn_tco229: string;
   attribute syn_tco229 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OUT = 2.966";
   attribute syn_tco230: string;
   attribute syn_tco230 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_H2F_A = 3.391";
   attribute syn_tco231: string;
   attribute syn_tco231 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_OUT = 3.117";
   attribute syn_tco232: string;
   attribute syn_tco232 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_A = 3.384";
   attribute syn_tco233: string;
   attribute syn_tco233 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_B = 3.436";
   attribute syn_tco234: string;
   attribute syn_tco234 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_OUT = 3.077";
   attribute syn_tco235: string;
   attribute syn_tco235 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_A = 3.508";
   attribute syn_tco236: string;
   attribute syn_tco236 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_B = 3.215";
   attribute syn_tco237: string;
   attribute syn_tco237 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_USBC_DATA3_MGPIO26B_OE = 3.090";
   attribute syn_tco238: string;
   attribute syn_tco238 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT = 3.048";
   attribute syn_tco239: string;
   attribute syn_tco239 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_A = 3.317";
   attribute syn_tco240: string;
   attribute syn_tco240 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_B = 3.509";
   attribute syn_tco241: string;
   attribute syn_tco241 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OE = 3.308";
   attribute syn_tco242: string;
   attribute syn_tco242 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT = 3.278";
   attribute syn_tco243: string;
   attribute syn_tco243 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_A = 3.464";
   attribute syn_tco244: string;
   attribute syn_tco244 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_B = 4.454";
   attribute syn_tco245: string;
   attribute syn_tco245 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OE = 3.467";
   attribute syn_tco246: string;
   attribute syn_tco246 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT = 3.318";
   attribute syn_tco247: string;
   attribute syn_tco247 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE = 3.954";
   attribute syn_tco248: string;
   attribute syn_tco248 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT = 4.201";
   attribute syn_tco249: string;
   attribute syn_tco249 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_A = 3.546";
   attribute syn_tco250: string;
   attribute syn_tco250 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_B = 3.547";
   attribute syn_tco251: string;
   attribute syn_tco251 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_A = 3.616";
   attribute syn_tco252: string;
   attribute syn_tco252 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_B = 3.530";
   attribute syn_tco253: string;
   attribute syn_tco253 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OUT = 5.270";
   attribute syn_tco254: string;
   attribute syn_tco254 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_A = 3.399";
   attribute syn_tco255: string;
   attribute syn_tco255 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_B = 3.503";
   attribute syn_tco256: string;
   attribute syn_tco256 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_A = 3.533";
   attribute syn_tco257: string;
   attribute syn_tco257 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_B = 3.558";
   attribute syn_tco258: string;
   attribute syn_tco258 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_USBA_DATA5_MGPIO8A_OE = 3.226";
   attribute syn_tco259: string;
   attribute syn_tco259 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_USBA_DATA5_MGPIO8A_OUT = 3.399";
   attribute syn_tco260: string;
   attribute syn_tco260 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_A = 3.368";
   attribute syn_tco261: string;
   attribute syn_tco261 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_B = 3.395";
   attribute syn_tco262: string;
   attribute syn_tco262 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_USBA_DATA6_MGPIO9A_OE = 3.132";
   attribute syn_tco263: string;
   attribute syn_tco263 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_USBA_DATA6_MGPIO9A_OUT = 3.275";
   attribute syn_tco264: string;
   attribute syn_tco264 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_A = 3.422";
   attribute syn_tco265: string;
   attribute syn_tco265 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_B = 3.482";
   attribute syn_tco266: string;
   attribute syn_tco266 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_USBA_DATA7_MGPIO10A_OE = 3.137";
   attribute syn_tco267: string;
   attribute syn_tco267 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_USBA_DATA7_MGPIO10A_OUT = 3.297";
   attribute syn_tco268: string;
   attribute syn_tco268 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS4_MGPIO19A_H2F_A = 3.563";
   attribute syn_tco269: string;
   attribute syn_tco269 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS5_MGPIO20A_H2F_A = 3.248";
   attribute syn_tco270: string;
   attribute syn_tco270 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS6_MGPIO21A_H2F_A = 3.435";
   attribute syn_tco271: string;
   attribute syn_tco271 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS7_MGPIO22A_H2F_A = 3.667";
   attribute syn_tco272: string;
   attribute syn_tco272 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_A = 3.621";
   attribute syn_tco273: string;
   attribute syn_tco273 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_B = 3.944";
   attribute syn_tco274: string;
   attribute syn_tco274 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_OE = 3.051";
   attribute syn_tco275: string;
   attribute syn_tco275 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_OUT = 3.503";
   attribute syn_tco276: string;
   attribute syn_tco276 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_A = 3.254";
   attribute syn_tco277: string;
   attribute syn_tco277 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_B = 3.406";
   attribute syn_tco278: string;
   attribute syn_tco278 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OE = 3.510";
   attribute syn_tco279: string;
   attribute syn_tco279 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OUT = 3.540";
   attribute syn_tco280: string;
   attribute syn_tco280 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_A = 3.869";
   attribute syn_tco281: string;
   attribute syn_tco281 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_B = 4.066";
   attribute syn_tco282: string;
   attribute syn_tco282 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_OE = 3.269";
   attribute syn_tco283: string;
   attribute syn_tco283 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_OUT = 3.379";
   attribute syn_tco284: string;
   attribute syn_tco284 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_A = 3.397";
   attribute syn_tco285: string;
   attribute syn_tco285 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_B = 3.268";
   attribute syn_tco286: string;
   attribute syn_tco286 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_OE = 3.393";
   attribute syn_tco287: string;
   attribute syn_tco287 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_OUT = 3.348";
   attribute syn_tco288: string;
   attribute syn_tco288 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_A = 3.442";
   attribute syn_tco289: string;
   attribute syn_tco289 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_B = 3.288";
   attribute syn_tco290: string;
   attribute syn_tco290 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_OE = 3.352";
   attribute syn_tco291: string;
   attribute syn_tco291 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_OUT = 3.195";
   attribute syn_tco292: string;
   attribute syn_tco292 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_A = 3.319";
   attribute syn_tco293: string;
   attribute syn_tco293 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_B = 3.381";
   attribute syn_tco294: string;
   attribute syn_tco294 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_OE = 3.460";
   attribute syn_tco295: string;
   attribute syn_tco295 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_OUT = 3.601";
   attribute syn_tco296: string;
   attribute syn_tco296 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_H2F_A = 3.689";
   attribute syn_tco297: string;
   attribute syn_tco297 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_OE = 3.404";
   attribute syn_tco298: string;
   attribute syn_tco298 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_OUT = 3.350";
   attribute syn_tco299: string;
   attribute syn_tco299 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_H2F_A = 3.385";
   attribute syn_tco300: string;
   attribute syn_tco300 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_OE = 3.501";
   attribute syn_tco301: string;
   attribute syn_tco301 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_OUT = 3.421";
   attribute syn_tco302: string;
   attribute syn_tco302 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_H2F_A = 3.501";
   attribute syn_tco303: string;
   attribute syn_tco303 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_OE = 3.267";
   attribute syn_tco304: string;
   attribute syn_tco304 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_OUT = 3.448";
   attribute syn_tco305: string;
   attribute syn_tco305 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_H2F_A = 3.443";
   attribute syn_tco306: string;
   attribute syn_tco306 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_OE = 3.380";
   attribute syn_tco307: string;
   attribute syn_tco307 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_OUT = 3.539";
   attribute black_box_pad_pin : string;
   attribute black_box_pad_pin of DEF_ARCH : architecture is "";

begin

end DEF_ARCH;
