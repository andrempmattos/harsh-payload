-- Version: v11.8 11.8.0.26

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity openbank is

    port( wshift_13               : out   std_logic_vector(6 downto 1);
          wshift                  : in    std_logic_vector(6 downto 1);
          raddr                   : in    std_logic_vector(22 downto 0);
          lnht_cmd                : in    std_logic_vector(3 downto 0);
          pcable                  : inout std_logic_vector(3 downto 0) := (others => 'Z');
          active                  : inout std_logic_vector(3 downto 0) := (others => 'Z');
          bdcnt                   : in    std_logic_vector(3 downto 0);
          rdwr_cmd                : in    std_logic_vector(3 downto 0);
          dorw                    : in    std_logic_vector(3 downto 0);
          rshift                  : in    std_logic_vector(6 downto 5);
          bcount                  : in    std_logic_vector(2 downto 0);
          line_i_2                : out   std_logic_vector(11 downto 0);
          bdcnt_6_iv_i_0          : out   std_logic;
          rwable_1                : in    std_logic;
          rwable_0                : in    std_logic;
          rwable_3                : in    std_logic;
          bdcnt_6_2               : out   std_logic;
          bdcnt_6_0               : out   std_logic;
          bdcnt_6_3               : out   std_logic;
          actable_2               : out   std_logic;
          actable_3               : in    std_logic;
          actable_0               : in    std_logic;
          cs_n_5_0                : out   std_logic;
          sa_5_5                  : out   std_logic;
          sa_5_1                  : out   std_logic;
          sa_5_0                  : out   std_logic;
          sa_5_10                 : out   std_logic;
          sa_5_8                  : out   std_logic;
          sa_5_2                  : out   std_logic;
          sa_5_3                  : out   std_logic;
          sa_5_4                  : out   std_logic;
          psa_0                   : in    std_logic;
          psa_8                   : in    std_logic;
          prch_0                  : in    std_logic;
          goact_2                 : in    std_logic;
          goact_0                 : in    std_logic;
          goact_3                 : in    std_logic;
          rshift_46_0             : out   std_logic;
          chip_i_2_0              : out   std_logic;
          rw_4                    : out   std_logic;
          N_117_i                 : out   std_logic;
          N_78_i                  : out   std_logic;
          un155_rdwr_cmd          : out   std_logic;
          un197_rdwr_cmd          : out   std_logic;
          un71_rdwr_cmd           : out   std_logic;
          un113_rdwr_cmd          : out   std_logic;
          pchaddr_3_sqmuxa_i_0    : out   std_logic;
          act_4                   : out   std_logic;
          un30_rdwr_cmd           : in    std_logic;
          un42_rdwr_cmd           : in    std_logic;
          N_783_i                 : out   std_logic;
          N_77                    : out   std_logic;
          oe_2                    : out   std_logic;
          w_valid_i               : in    std_logic;
          rc_zero_0_sqmuxa        : out   std_logic;
          wc_zero_0_sqmuxa        : out   std_logic;
          N_812                   : in    std_logic;
          un222_rdwr_cmd          : out   std_logic;
          un180_rdwr_cmd          : out   std_logic;
          un18_rdwr_cmd           : out   std_logic;
          un54_rdwr_cmd           : out   std_logic;
          un138_rdwr_cmd          : out   std_logic;
          un7_mode_cmd            : out   std_logic;
          un13_rfsh_cmd           : out   std_logic;
          N_73                    : in    std_logic;
          un13_rfsh_cmd_1         : in    std_logic;
          we_n_2                  : out   std_logic;
          un16_act_i              : in    std_logic;
          un1_pch_3_i             : out   std_logic;
          un96_rdwr_cmd           : out   std_logic;
          un1_cs_n_0_sqmuxa_i_0   : in    std_logic;
          bdzero_2                : out   std_logic;
          bterm_3                 : out   std_logic;
          w_valid_i_1             : out   std_logic;
          rcount_2_sqmuxa         : out   std_logic;
          un217_rdwr_cmd          : out   std_logic;
          turnaround_hold         : in    std_logic;
          rc_zero_d               : in    std_logic;
          un1_mode_cmd            : out   std_logic;
          mode_cmd                : in    std_logic;
          refresh                 : in    std_logic;
          un4_p_req_0_49_a2_0_a2  : out   std_logic;
          p_req                   : in    std_logic;
          un1_pch_4_1             : out   std_logic;
          bterm                   : in    std_logic;
          pchaddr_9_sn_m2_i_1     : out   std_logic;
          pchaddr_9_sn_m3_i_1     : out   std_logic;
          mode                    : in    std_logic;
          read_cmd                : in    std_logic;
          un4_rf_req_0_60_a2_0_a2 : out   std_logic;
          rf_req                  : in    std_logic;
          precharge               : in    std_logic;
          doread                  : in    std_logic;
          un36_rw_i_0             : out   std_logic;
          un13_prch_cmd           : out   std_logic;
          rfsh_cmd                : in    std_logic;
          prch_cmd                : in    std_logic;
          bdzero                  : in    std_logic;
          un14_rw                 : in    std_logic;
          N_125                   : out   std_logic;
          bterm_cmd               : in    std_logic;
          ack                     : in    std_logic;
          lnht_cmd26              : out   std_logic;
          un1_rowaddr_int_0_N_2   : in    std_logic;
          lnht_cmd5               : out   std_logic;
          un1_line_i_0_0_N_2      : in    std_logic;
          cke                     : in    std_logic;
          un8_rc_zero             : out   std_logic;
          rc_zero                 : in    std_logic;
          un4_wc_zero             : out   std_logic;
          wc_zero                 : in    std_logic;
          dowrite                 : in    std_logic;
          rw                      : in    std_logic;
          sa_5_sn_N_4_mux         : in    std_logic;
          N_6                     : in    std_logic;
          un78_rw                 : in    std_logic;
          un1_rw_11_i             : out   std_logic;
          pch                     : in    std_logic;
          un8_precharge           : in    std_logic;
          act                     : in    std_logic;
          clk                     : in    std_logic;
          reset_n                 : in    std_logic
        );

end openbank;

architecture DEF_ARCH of openbank is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \actable_shift[8]_net_1\, GND_net_1, 
        \actable_shift_57[8]_net_1\, VCC_net_1, 
        \actable_shift[9]_net_1\, \actable_shift_57[9]_net_1\, 
        \actable_shift[10]_net_1\, \actable_shift_57[10]_net_1\, 
        \actable_shift[11]_net_1\, \actable_shift_57[11]_net_1\, 
        \actable_shift[12]_net_1\, \actable_shift_57[12]_net_1\, 
        \pcable_shift[3]_net_1\, N_752_i, \pcable_shift[4]_net_1\, 
        \pcable_shift_13[4]\, \pcable_shift[5]_net_1\, 
        \pcable_shift_13[5]\, \pcable_shift[6]_net_1\, N_4_i, 
        \pcable_shift[7]_net_1\, \pcable_shift_13[7]\, 
        \pcable_shift[8]_net_1\, \pcable_shift_0_sqmuxa_i\, 
        \rc_shift[7]_net_1\, \rc_shift_30[7]_net_1\, 
        \rwable_shift[0]_net_1\, \rwable_shift_7[0]\, 
        \rwable_shift[1]_net_1\, \rwable_shift_7[1]\, 
        \rwable_shift[2]_net_1\, \rwable_shift_7[2]\, 
        \rwable_shift[3]_net_1\, \rwable_shift_7[3]\, 
        \rwable_shift[4]_net_1\, \rwable_shift_7[4]\, 
        \actable_shift[0]_net_1\, \actable_shift_57[0]_net_1\, 
        \actable_shift[1]_net_1\, \actable_shift_57[1]_net_1\, 
        \actable_shift[2]_net_1\, \actable_shift_57[2]_net_1\, 
        \actable_shift[3]_net_1\, \actable_shift_57[3]_net_1\, 
        \actable_shift[4]_net_1\, \actable_shift_57[4]_net_1\, 
        \actable_shift[5]_net_1\, \actable_shift_57[5]_net_1\, 
        \actable_shift[6]_net_1\, \actable_shift_57[6]_net_1\, 
        \actable_shift[7]_net_1\, \actable_shift_57[7]_net_1\, 
        \rc_shift[0]_net_1\, \rc_shift_30[0]_net_1\, 
        \rc_shift[1]_net_1\, \rc_shift_30[1]_net_1\, 
        \rc_shift[2]_net_1\, \rc_shift_30[2]_net_1\, 
        \rc_shift[3]_net_1\, \rc_shift_30[3]_net_1\, 
        \rc_shift[4]_net_1\, \rc_shift_30[4]_net_1\, 
        \rc_shift[5]_net_1\, \rc_shift_30[5]_net_1\, 
        \rc_shift[6]_net_1\, \rc_shift_30[6]_net_1\, un36_dopch, 
        \prev_cmd_read\, \prev_cmd_read_1\, N_751_i, \rwable[2]\, 
        rwable_int_3, actable_6, N_331_i, sa_5_0_0, sa_5, 
        \rshift_46_1[5]\, \un1_rw_11_i\, \sa_5_1[5]\, \sa_5_1[1]\, 
        \sa_5_1[0]\, un197_rdwr_cmd_0_a2_1, un71_rdwr_cmd_0_a2_1, 
        rw_4_0_a2_1, un113_rdwr_cmd_0_a2_1, N_756, un47_rw, 
        un5_dopch_i, \N_125\, \CO1\, bdzero_0_sqmuxa, un4_bdzero, 
        \un36_rw_i_0\, doread_m, N_68, \un1_goactive_4_1\, 
        un96_rdwr_cmd_0_a2_2, un180_rdwr_cmd_0_a2_1, 
        un138_rdwr_cmd_0_a2_1, un36_rw_i_0_3, N_126, un9_bdzero, 
        N_122, \actable_1_sqmuxa_2\, \un217_rdwr_cmd\, un20_rw, 
        un28_rw, \w_valid_i_1\, bdcnt_2_sqmuxa, 
        \bdcnt_6_iv_0_0[1]\, \un96_rdwr_cmd\, \un1_pch_3_i\, 
        \un138_rdwr_cmd\, \un54_rdwr_cmd\, \un18_rdwr_cmd\, 
        un1_goactive_4_i, \un180_rdwr_cmd\, \un222_rdwr_cmd\, 
        actable_shift_57_sm0, N_130, \actable_shift_57_ss0\, 
        \actable_shift_57_m2[12]_net_1\, 
        \actable_shift_57_m2[11]_net_1\, 
        \actable_shift_57_m2[10]_net_1\, 
        \actable_shift_57_m2[9]_net_1\, 
        \actable_shift_57_m2[8]_net_1\, 
        \actable_shift_57_m2[7]_net_1\, 
        \actable_shift_57_m2[6]_net_1\, 
        \actable_shift_57_m2[5]_net_1\, 
        \actable_shift_57_m2[4]_net_1\, 
        \actable_shift_57_m2[3]_net_1\, 
        \actable_shift_57_m2[2]_net_1\, 
        \actable_shift_57_m2[1]_net_1\, \un113_rdwr_cmd\, 
        \un71_rdwr_cmd\, \un197_rdwr_cmd\, \un155_rdwr_cmd\
         : std_logic;

begin 

    un155_rdwr_cmd <= \un155_rdwr_cmd\;
    un197_rdwr_cmd <= \un197_rdwr_cmd\;
    un71_rdwr_cmd <= \un71_rdwr_cmd\;
    un113_rdwr_cmd <= \un113_rdwr_cmd\;
    un222_rdwr_cmd <= \un222_rdwr_cmd\;
    un180_rdwr_cmd <= \un180_rdwr_cmd\;
    un18_rdwr_cmd <= \un18_rdwr_cmd\;
    un54_rdwr_cmd <= \un54_rdwr_cmd\;
    un138_rdwr_cmd <= \un138_rdwr_cmd\;
    un1_pch_3_i <= \un1_pch_3_i\;
    un96_rdwr_cmd <= \un96_rdwr_cmd\;
    w_valid_i_1 <= \w_valid_i_1\;
    un217_rdwr_cmd <= \un217_rdwr_cmd\;
    un36_rw_i_0 <= \un36_rw_i_0\;
    N_125 <= \N_125\;
    un1_rw_11_i <= \un1_rw_11_i\;

    \sd_ctl_p.sa_5_0\ : CFG4
      generic map(INIT => x"A080")

      port map(A => act, B => un8_precharge, C => psa_0, D => pch, 
        Y => sa_5_0_0);
    
    \line[4]\ : SLE
      port map(D => raddr(14), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(4));
    
    \rw_p.rwable_shift_7[3]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_2, B => un5_dopch_i, C => 
        \rwable_shift[4]_net_1\, Y => \rwable_shift_7[3]\);
    
    \actable_shift_57[9]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[9]_net_1\, C => 
        \actable_shift[10]_net_1\, D => refresh, Y => 
        \actable_shift_57[9]_net_1\);
    
    \line[1]\ : SLE
      port map(D => raddr(11), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(1));
    
    \pcable_shift[5]\ : SLE
      port map(D => \pcable_shift_13[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[5]_net_1\);
    
    \actable_shift[6]\ : SLE
      port map(D => \actable_shift_57[6]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[6]_net_1\);
    
    \rc_shift[6]\ : SLE
      port map(D => \rc_shift_30[6]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[6]_net_1\);
    
    \actable_shift_57_m2[10]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[11]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[10]_net_1\);
    
    \act_p.0.un71_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => rwable_0, B => lnht_cmd(0), C => 
        un71_rdwr_cmd_0_a2_1, D => N_130, Y => \un71_rdwr_cmd\);
    
    \sd_ctl_p.we_n_2_iv_RNO\ : CFG2
      generic map(INIT => x"8")

      port map(A => \un36_rw_i_0\, B => doread, Y => doread_m);
    
    \act_p.1.un113_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => rwable_1, B => lnht_cmd(1), C => 
        un113_rdwr_cmd_0_a2_1, D => N_130, Y => \un113_rdwr_cmd\);
    
    \actable_shift_57_m2[1]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[2]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[1]_net_1\);
    
    \line[8]\ : SLE
      port map(D => raddr(18), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(8));
    
    \bterm_p.op_eq.un9_bdzero_RNIDJGS\ : CFG4
      generic map(INIT => x"00E4")

      port map(A => rw, B => un9_bdzero, C => un28_rw, D => N_68, 
        Y => N_783_i);
    
    \sd_ctl_p.sa_5\ : CFG4
      generic map(INIT => x"5040")

      port map(A => act, B => un8_precharge, C => psa_0, D => pch, 
        Y => sa_5);
    
    \rc_shift[1]\ : SLE
      port map(D => \rc_shift_30[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[1]_net_1\);
    
    \pcable_shift_RNO[7]\ : CFG4
      generic map(INIT => x"2AAA")

      port map(A => \pcable_shift[8]_net_1\, B => dorw(2), C => 
        bcount(1), D => bcount(2), Y => \pcable_shift_13[7]\);
    
    \actable_shift_57_m2[9]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[10]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[9]_net_1\);
    
    un5_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => precharge, B => prch_0, Y => un5_dopch_i);
    
    \actable_shift_57[8]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[8]_net_1\, C => 
        \actable_shift[9]_net_1\, D => refresh, Y => 
        \actable_shift_57[8]_net_1\);
    
    \line[9]\ : SLE
      port map(D => raddr(19), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(9));
    
    \bterm_p.bdcnt_6_iv_i[1]\ : CFG4
      generic map(INIT => x"3233")

      port map(A => un28_rw, B => \bdcnt_6_iv_0_0[1]\, C => 
        bcount(1), D => rw, Y => bdcnt_6_iv_i_0);
    
    \actable_shift[12]\ : SLE
      port map(D => \actable_shift_57[12]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[12]_net_1\);
    
    un1_goactive_4 : CFG3
      generic map(INIT => x"10")

      port map(A => refresh, B => un5_dopch_i, C => 
        \un1_goactive_4_1\, Y => un1_goactive_4_i);
    
    \line[3]\ : SLE
      port map(D => raddr(13), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(3));
    
    \sd_ctl_p.sa_5[4]\ : CFG4
      generic map(INIT => x"C840")

      port map(A => act, B => sa_5_sn_N_4_mux, C => raddr(4), D
         => raddr(14), Y => sa_5_4);
    
    \act_p.rw_4_0_a2_1\ : CFG4
      generic map(INIT => x"B000")

      port map(A => rc_zero_d, B => turnaround_hold, C => 
        read_cmd, D => rc_zero, Y => N_122);
    
    pcable_int : SLE
      port map(D => N_751_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => pcable(2));
    
    \actable_shift_57[3]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[3]_net_1\, Y => 
        \actable_shift_57[3]_net_1\);
    
    \rc_shift[3]\ : SLE
      port map(D => \rc_shift_30[3]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[3]_net_1\);
    
    \act_p.3.un217_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(3), B => active(3), C => pcable(3), 
        D => lnht_cmd(3), Y => \un217_rdwr_cmd\);
    
    \act_p.1.un138_rdwr_cmd_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => un138_rdwr_cmd_0_a2_1, B => bterm_cmd, C => 
        pch, Y => \un138_rdwr_cmd\);
    
    \dh_p.un35_mode_cmd_i_a2\ : CFG3
      generic map(INIT => x"01")

      port map(A => prch_cmd, B => mode_cmd, C => rfsh_cmd, Y => 
        N_126);
    
    \act_p.rw_4_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \rwable[2]\, B => lnht_cmd(2), C => 
        rw_4_0_a2_1, D => N_130, Y => \un155_rdwr_cmd\);
    
    \rc_zero_0_sqmuxa\ : CFG2
      generic map(INIT => x"8")

      port map(A => un78_rw, B => N_812, Y => rc_zero_0_sqmuxa);
    
    \cmd_p.3.lnht_cmd26\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_rowaddr_int_0_N_2, B => goact_3, Y => 
        lnht_cmd26);
    
    un7_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => un5_dopch_i, B => goact_2, Y => un36_dopch);
    
    \cmd_p.0.lnht_cmd5\ : CFG2
      generic map(INIT => x"D")

      port map(A => un1_line_i_0_0_N_2, B => goact_0, Y => 
        lnht_cmd5);
    
    pcable_int_RNISSEN : CFG4
      generic map(INIT => x"FF7F")

      port map(A => rdwr_cmd(2), B => active(2), C => pcable(2), 
        D => lnht_cmd(2), Y => pchaddr_9_sn_m2_i_1);
    
    \actable_shift_57[10]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[10]_net_1\, C => 
        \actable_shift[11]_net_1\, D => refresh, Y => 
        \actable_shift_57[10]_net_1\);
    
    \rc_shift_30[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_2, B => \rc_shift[6]_net_1\, Y => 
        \rc_shift_30[5]_net_1\);
    
    \line[5]\ : SLE
      port map(D => raddr(15), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(5));
    
    pcable_int_RNO : CFG4
      generic map(INIT => x"0E04")

      port map(A => \prev_cmd_read\, B => \pcable_shift[3]_net_1\, 
        C => dorw(2), D => \pcable_shift[4]_net_1\, Y => N_751_i);
    
    \actable_shift[8]\ : SLE
      port map(D => \actable_shift_57[8]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[8]_net_1\);
    
    \pcable_shift[6]\ : SLE
      port map(D => N_4_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[6]_net_1\);
    
    \act_p.rw_4_0_a2_0\ : CFG4
      generic map(INIT => x"F040")

      port map(A => read_cmd, B => wc_zero, C => \N_125\, D => 
        N_122, Y => N_130);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \act_p.0.un18_rdwr_cmd_0_a2_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => ack, B => bterm_cmd, Y => \N_125\);
    
    \actable_shift_57_m2[12]\ : CFG3
      generic map(INIT => x"54")

      port map(A => active(2), B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_m2[12]_net_1\);
    
    \sd_ctl_p.cs_n_5_0_a2[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => mode, B => precharge, C => 
        un1_cs_n_0_sqmuxa_i_0, D => refresh, Y => cs_n_5_0);
    
    \psa_p.un13_prch_cmd\ : CFG2
      generic map(INIT => x"E")

      port map(A => prch_cmd, B => rfsh_cmd, Y => un13_prch_cmd);
    
    \rc_shift_30[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_2, B => \rc_shift[1]_net_1\, Y => 
        \rc_shift_30[0]_net_1\);
    
    \act_p.pchaddr_9_sn_m3_i_1\ : CFG4
      generic map(INIT => x"FF7F")

      port map(A => rdwr_cmd(1), B => active(1), C => pcable(1), 
        D => lnht_cmd(1), Y => pchaddr_9_sn_m3_i_1);
    
    actable_1_sqmuxa_2 : CFG4
      generic map(INIT => x"0008")

      port map(A => \rc_shift[0]_net_1\, B => mode, C => refresh, 
        D => un5_dopch_i, Y => \actable_1_sqmuxa_2\);
    
    \sd_ctl_p.sa_5[0]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => sa_5, B => sa_5_sn_N_4_mux, C => \sa_5_1[0]\, 
        D => sa_5_0_0, Y => sa_5_0);
    
    \act_p.0.un71_rdwr_cmd_0_a2_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => dorw(0), B => rdwr_cmd(0), Y => 
        un71_rdwr_cmd_0_a2_1);
    
    \sd_ctl_p.sa_5[10]\ : CFG4
      generic map(INIT => x"B830")

      port map(A => act, B => sa_5_sn_N_4_mux, C => psa_8, D => 
        raddr(20), Y => sa_5_10);
    
    \line[11]\ : SLE
      port map(D => raddr(21), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(11));
    
    \bterm_p.bdcnt_6_iv_0_0[1]\ : CFG4
      generic map(INIT => x"CEEC")

      port map(A => un4_bdzero, B => N_68, C => bdcnt(1), D => 
        bdcnt(0), Y => \bdcnt_6_iv_0_0[1]\);
    
    \actable_shift_57_m2[5]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[6]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[5]_net_1\);
    
    \line[10]\ : SLE
      port map(D => raddr(20), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(10));
    
    prev_cmd_read : SLE
      port map(D => \prev_cmd_read_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \prev_cmd_read\);
    
    \actable_shift[10]\ : SLE
      port map(D => \actable_shift_57[10]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[10]_net_1\);
    
    \pcable_shift_RNO[6]\ : CFG4
      generic map(INIT => x"02AA")

      port map(A => \pcable_shift[7]_net_1\, B => bcount(0), C
         => bcount(1), D => N_756, Y => N_4_i);
    
    \act_p.un13_rfsh_cmd_0_a2\ : CFG3
      generic map(INIT => x"04")

      port map(A => refresh, B => un13_rfsh_cmd_1, C => N_73, Y
         => un13_rfsh_cmd);
    
    \act_p.act_4_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un54_rdwr_cmd\, B => un42_rdwr_cmd, C => 
        un30_rdwr_cmd, D => \un18_rdwr_cmd\, Y => act_4);
    
    \cmd_p.un4_rf_req_0_60_a2_0_a2\ : CFG2
      generic map(INIT => x"4")

      port map(A => ack, B => rf_req, Y => 
        un4_rf_req_0_60_a2_0_a2);
    
    \dh_p.un35_mode_cmd_i_a2_RNIRT47\ : CFG3
      generic map(INIT => x"01")

      port map(A => ack, B => N_126, C => N_73, Y => N_78_i);
    
    \act_p.rw_4_0_a2_1_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => dorw(2), B => rdwr_cmd(2), Y => rw_4_0_a2_1);
    
    \actable_shift_57[11]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[11]_net_1\, C => 
        \actable_shift[12]_net_1\, D => refresh, Y => 
        \actable_shift_57[11]_net_1\);
    
    \wshift_13[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => un47_rw, B => wshift(4), C => bcount(2), Y
         => wshift_13(3));
    
    \actable_shift_57[2]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[2]_net_1\, Y => 
        \actable_shift_57[2]_net_1\);
    
    un36_rw : CFG2
      generic map(INIT => x"8")

      port map(A => un36_rw_i_0_3, B => rw, Y => \un36_rw_i_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \rc_shift[4]\ : SLE
      port map(D => \rc_shift_30[4]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[4]_net_1\);
    
    \rc_p.un8_rc_zero_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => rw, B => rc_zero, Y => un8_rc_zero);
    
    \bterm_p.bdcnt_6_0_iv[2]\ : CFG4
      generic map(INIT => x"BA30")

      port map(A => bcount(2), B => N_331_i, C => un4_bdzero, D
         => bdcnt_2_sqmuxa, Y => bdcnt_6_2);
    
    \actable_shift[5]\ : SLE
      port map(D => \actable_shift_57[5]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[5]_net_1\);
    
    \rcount_2_sqmuxa\ : CFG2
      generic map(INIT => x"8")

      port map(A => un47_rw, B => bcount(2), Y => rcount_2_sqmuxa);
    
    \actable_shift_57[0]\ : CFG4
      generic map(INIT => x"00EA")

      port map(A => un5_dopch_i, B => \actable_shift_57_ss0\, C
         => \actable_shift[1]_net_1\, D => refresh, Y => 
        \actable_shift_57[0]_net_1\);
    
    \pcable_shift[3]\ : SLE
      port map(D => N_752_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[3]_net_1\);
    
    \actable_shift_57[6]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[6]_net_1\, C => 
        \actable_shift[7]_net_1\, D => refresh, Y => 
        \actable_shift_57[6]_net_1\);
    
    prev_cmd_read_1 : CFG3
      generic map(INIT => x"D8")

      port map(A => dorw(2), B => read_cmd, C => \prev_cmd_read\, 
        Y => \prev_cmd_read_1\);
    
    \pcable_shift_RNO[5]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[6]_net_1\, B => dorw(2), C => 
        bcount(2), Y => \pcable_shift_13[5]\);
    
    \actable_shift_57_m2[11]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[12]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[11]_net_1\);
    
    un1_rw_11_RNI72UI1 : CFG4
      generic map(INIT => x"E255")

      port map(A => \rshift_46_1[5]\, B => \un1_rw_11_i\, C => 
        rshift(5), D => un78_rw, Y => rshift_46_0);
    
    \rwable_shift[2]\ : SLE
      port map(D => \rwable_shift_7[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[2]_net_1\);
    
    \actable_shift_57_m2[7]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[8]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[7]_net_1\);
    
    \wc_p.un47_rw\ : CFG2
      generic map(INIT => x"8")

      port map(A => rw, B => dowrite, Y => un47_rw);
    
    \act_p.un7_mode_cmd\ : CFG3
      generic map(INIT => x"02")

      port map(A => mode_cmd, B => mode, C => N_73, Y => 
        un7_mode_cmd);
    
    \sd_ctl_p.sa_5_1[0]\ : CFG3
      generic map(INIT => x"47")

      port map(A => raddr(10), B => act, C => raddr(0), Y => 
        \sa_5_1[0]\);
    
    \cmd_p.un4_p_req_0_49_a2_0_a2\ : CFG3
      generic map(INIT => x"04")

      port map(A => rf_req, B => p_req, C => ack, Y => 
        un4_p_req_0_49_a2_0_a2);
    
    \bterm_p.op_eq.un9_bdzero\ : CFG4
      generic map(INIT => x"1000")

      port map(A => bdcnt(3), B => bdcnt(2), C => bdcnt(1), D => 
        bdcnt(0), Y => un9_bdzero);
    
    \bterm_p.bterm_3_iv\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un4_bdzero, B => bdzero_0_sqmuxa, C => 
        bterm_cmd, Y => bterm_3);
    
    un1_goactive_4_1 : CFG4
      generic map(INIT => x"0031")

      port map(A => act, B => goact_2, C => active(2), D => mode, 
        Y => \un1_goactive_4_1\);
    
    \actable_shift_57_m2[6]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[7]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[6]_net_1\);
    
    \rc_shift_30[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_2, B => cke, Y => 
        \rc_shift_30[7]_net_1\);
    
    \actable_shift_57_m2[2]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[3]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[2]_net_1\);
    
    \wshift_13[5]\ : CFG4
      generic map(INIT => x"B830")

      port map(A => bcount(2), B => un47_rw, C => wshift(6), D
         => bcount(1), Y => wshift_13(5));
    
    \act_p.0.un96_rdwr_cmd_0_a2_2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(0), B => active(0), C => pcable(0), 
        D => lnht_cmd(0), Y => un96_rdwr_cmd_0_a2_2);
    
    \wshift_13[6]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => bcount(0), B => bcount(1), C => bcount(2), D
         => un47_rw, Y => wshift_13(6));
    
    \wshift_13[1]\ : CFG3
      generic map(INIT => x"4E")

      port map(A => un47_rw, B => wshift(2), C => un20_rw, Y => 
        wshift_13(1));
    
    \act_p.2.un180_rdwr_cmd_0_a2_1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(2), B => active(2), C => pcable(2), 
        D => lnht_cmd(2), Y => un180_rdwr_cmd_0_a2_1);
    
    \actable_shift_57_m2[3]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[4]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[3]_net_1\);
    
    \rw_p.rwable_shift_7[4]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => active(2), B => goact_2, C => un5_dopch_i, Y
         => \rwable_shift_7[4]\);
    
    \actable_shift_57[5]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[5]_net_1\, Y => 
        \actable_shift_57[5]_net_1\);
    
    \actable_shift[4]\ : SLE
      port map(D => \actable_shift_57[4]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[4]_net_1\);
    
    \wshift_13[2]\ : CFG4
      generic map(INIT => x"3074")

      port map(A => un28_rw, B => un47_rw, C => wshift(3), D => 
        un20_rw, Y => wshift_13(2));
    
    \un1_pch_4_1\ : CFG3
      generic map(INIT => x"04")

      port map(A => bterm, B => pch, C => rw, Y => un1_pch_4_1);
    
    \rc_shift[2]\ : SLE
      port map(D => \rc_shift_30[2]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[2]_net_1\);
    
    \line[0]\ : SLE
      port map(D => raddr(10), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(0));
    
    \rw_p.rwable_shift_7[2]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_2, B => un5_dopch_i, C => 
        \rwable_shift[3]_net_1\, Y => \rwable_shift_7[2]\);
    
    \pcable_shift[7]\ : SLE
      port map(D => \pcable_shift_13[7]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[7]_net_1\);
    
    \bterm_p.op_eq.un20_rw\ : CFG3
      generic map(INIT => x"02")

      port map(A => bcount(0), B => bcount(1), C => bcount(2), Y
         => un20_rw);
    
    \rw_p.rwable_int_3_iv\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_2, B => un5_dopch_i, C => 
        \rwable_shift[0]_net_1\, Y => rwable_int_3);
    
    \act_p.1.un138_rdwr_cmd_0_a2_1\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(1), B => active(1), C => pcable(1), 
        D => lnht_cmd(1), Y => un138_rdwr_cmd_0_a2_1);
    
    \act_p.3.un197_rdwr_cmd_0_a2_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => dorw(3), B => rdwr_cmd(3), Y => 
        un197_rdwr_cmd_0_a2_1);
    
    \rc_shift[7]\ : SLE
      port map(D => \rc_shift_30[7]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[7]_net_1\);
    
    \act_p.2.un180_rdwr_cmd_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => un180_rdwr_cmd_0_a2_1, B => bterm_cmd, C => 
        pch, Y => \un180_rdwr_cmd\);
    
    \act_p.rw_4_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un197_rdwr_cmd\, B => \un155_rdwr_cmd\, C
         => \un113_rdwr_cmd\, D => \un71_rdwr_cmd\, Y => rw_4);
    
    \rc_shift_30[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_2, B => \rc_shift[4]_net_1\, Y => 
        \rc_shift_30[3]_net_1\);
    
    \line[7]\ : SLE
      port map(D => raddr(17), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(7));
    
    rwable_int : SLE
      port map(D => rwable_int_3, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rwable[2]\);
    
    \actable_shift[3]\ : SLE
      port map(D => \actable_shift_57[3]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[3]_net_1\);
    
    \act_p.0.un96_rdwr_cmd_0_a2\ : CFG3
      generic map(INIT => x"02")

      port map(A => un96_rdwr_cmd_0_a2_2, B => bterm_cmd, C => 
        pch, Y => \un96_rdwr_cmd\);
    
    \rc_shift_30[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_2, B => \rc_shift[7]_net_1\, Y => 
        \rc_shift_30[6]_net_1\);
    
    \sd_ctl_p.we_n_2_iv\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un16_act_i, B => refresh, C => doread_m, D
         => \un1_pch_3_i\, Y => we_n_2);
    
    \rc_shift[0]\ : SLE
      port map(D => \rc_shift_30[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[0]_net_1\);
    
    \actable_shift[1]\ : SLE
      port map(D => \actable_shift_57[1]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[1]_net_1\);
    
    \bterm_p.un4_bdzero_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => rw, B => bdzero, Y => un4_bdzero);
    
    pcable_shift_0_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bcount(1), B => bcount(2), C => dorw(2), D
         => bcount(0), Y => \pcable_shift_0_sqmuxa_i\);
    
    \actable_shift_57[4]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[4]_net_1\, Y => 
        \actable_shift_57[4]_net_1\);
    
    \pcable_shift[4]\ : SLE
      port map(D => \pcable_shift_13[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[4]_net_1\);
    
    \wr_flow_ctrl_p.oe_2\ : CFG2
      generic map(INIT => x"E")

      port map(A => \w_valid_i_1\, B => w_valid_i, Y => oe_2);
    
    \wc_zero_0_sqmuxa\ : CFG2
      generic map(INIT => x"8")

      port map(A => un47_rw, B => N_812, Y => wc_zero_0_sqmuxa);
    
    \rw_p.rwable_shift_7[0]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_2, B => un5_dopch_i, C => 
        \rwable_shift[1]_net_1\, Y => \rwable_shift_7[0]\);
    
    active_int : SLE
      port map(D => goact_2, CLK => clk, EN => un36_dopch, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => active(2));
    
    \actable_shift_57[7]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[7]_net_1\, C => 
        \actable_shift[8]_net_1\, D => refresh, Y => 
        \actable_shift_57[7]_net_1\);
    
    \sd_ctl_p.sa_5[5]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => sa_5, B => sa_5_sn_N_4_mux, C => \sa_5_1[5]\, 
        D => sa_5_0_0, Y => sa_5_5);
    
    bdzero_0_sqmuxa_0_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => un14_rw, B => rw, Y => bdzero_0_sqmuxa);
    
    \act_p.3.un217_rdwr_cmd_0_a2_RNI89HJ_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => pch, B => \un217_rdwr_cmd\, C => bterm_cmd, Y
         => \un222_rdwr_cmd\);
    
    \wc_p.un4_wc_zero_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => rw, B => wc_zero, Y => un4_wc_zero);
    
    \sd_ctl_p.sa_5_1[5]\ : CFG3
      generic map(INIT => x"47")

      port map(A => raddr(15), B => act, C => raddr(5), Y => 
        \sa_5_1[5]\);
    
    \data_flow_ctrl_p.rshift_46_1[5]\ : CFG3
      generic map(INIT => x"47")

      port map(A => N_6, B => un78_rw, C => rshift(6), Y => 
        \rshift_46_1[5]\);
    
    \pcable_shift[8]\ : SLE
      port map(D => \pcable_shift_0_sqmuxa_i\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[8]_net_1\);
    
    \actable_shift_57_m2[8]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[9]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[8]_net_1\);
    
    \wr_flow_ctrl_p.w_valid_i_1\ : CFG2
      generic map(INIT => x"E")

      port map(A => un47_rw, B => wshift(1), Y => \w_valid_i_1\);
    
    \rc_shift_30[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_2, B => \rc_shift[3]_net_1\, Y => 
        \rc_shift_30[2]_net_1\);
    
    \wshift_13[4]\ : CFG3
      generic map(INIT => x"4E")

      port map(A => un47_rw, B => wshift(5), C => N_6, Y => 
        wshift_13(4));
    
    \bterm_p.bdcnt_6_0_iv_RNO[2]\ : CFG3
      generic map(INIT => x"56")

      port map(A => bdcnt(2), B => bdcnt(1), C => bdcnt(0), Y => 
        N_331_i);
    
    \sd_ctl_p.sa_5[8]\ : CFG4
      generic map(INIT => x"B830")

      port map(A => act, B => sa_5_sn_N_4_mux, C => psa_8, D => 
        raddr(18), Y => sa_5_8);
    
    \line[6]\ : SLE
      port map(D => raddr(16), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(6));
    
    \bterm_p.bdzero_2_iv_0\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un4_bdzero, B => N_68, C => bterm_cmd, Y => 
        bdzero_2);
    
    \rwable_shift[3]\ : SLE
      port map(D => \rwable_shift_7[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[3]_net_1\);
    
    \actable_shift[0]\ : SLE
      port map(D => \actable_shift_57[0]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[0]_net_1\);
    
    un36_rw_3 : CFG4
      generic map(INIT => x"0001")

      port map(A => act, B => refresh, C => precharge, D => mode, 
        Y => un36_rw_i_0_3);
    
    \dh_p.un35_mode_cmd_i_a2_RNI4N87\ : CFG4
      generic map(INIT => x"AAAB")

      port map(A => rw, B => ack, C => N_73, D => N_126, Y => 
        N_117_i);
    
    actable_shift_57_m2s2 : CFG4
      generic map(INIT => x"FF02")

      port map(A => act, B => goact_2, C => active(2), D => mode, 
        Y => actable_shift_57_sm0);
    
    \pchaddr_3_sqmuxa_i_0\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un96_rdwr_cmd\, B => \un180_rdwr_cmd\, C => 
        \un138_rdwr_cmd\, D => \un222_rdwr_cmd\, Y => 
        pchaddr_3_sqmuxa_i_0);
    
    \actable_shift[9]\ : SLE
      port map(D => \actable_shift_57[9]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[9]_net_1\);
    
    \actable_shift_57[1]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[1]_net_1\, Y => 
        \actable_shift_57[1]_net_1\);
    
    \bterm_p.bdcnt_6_0_iv[0]\ : CFG4
      generic map(INIT => x"DC50")

      port map(A => bdcnt(0), B => bcount(0), C => un4_bdzero, D
         => bdcnt_2_sqmuxa, Y => bdcnt_6_0);
    
    \bterm_p.op_eq.un28_rw\ : CFG3
      generic map(INIT => x"04")

      port map(A => bcount(0), B => bcount(1), C => bcount(2), Y
         => un28_rw);
    
    bdcnt_2_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"04")

      port map(A => un28_rw, B => rw, C => un14_rw, Y => 
        bdcnt_2_sqmuxa);
    
    \act_p.3.un54_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(3), B => actable_3, C => \N_125\, D
         => goact_3, Y => \un54_rdwr_cmd\);
    
    un1_pcable_shift_3_sqmuxa_i_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => bcount(2), B => dorw(2), Y => N_756);
    
    \act_p.0.un18_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => rdwr_cmd(0), B => actable_0, C => \N_125\, D
         => goact_0, Y => \un18_rdwr_cmd\);
    
    \rw_p.rwable_shift_7[1]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_2, B => un5_dopch_i, C => 
        \rwable_shift[2]_net_1\, Y => \rwable_shift_7[1]\);
    
    \chip[0]\ : SLE
      port map(D => raddr(22), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => chip_i_2_0);
    
    \line[2]\ : SLE
      port map(D => raddr(12), CLK => clk, EN => goact_2, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_2(2));
    
    \sd_ctl_p.sa_5[1]\ : CFG4
      generic map(INIT => x"FFAE")

      port map(A => sa_5, B => sa_5_sn_N_4_mux, C => \sa_5_1[1]\, 
        D => sa_5_0_0, Y => sa_5_1);
    
    \actable_shift[11]\ : SLE
      port map(D => \actable_shift_57[11]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[11]_net_1\);
    
    \rwable_shift[0]\ : SLE
      port map(D => \rwable_shift_7[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[0]_net_1\);
    
    \rc_shift[5]\ : SLE
      port map(D => \rc_shift_30[5]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[5]_net_1\);
    
    \rwable_shift[1]\ : SLE
      port map(D => \rwable_shift_7[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[1]_net_1\);
    
    \rc_shift_30[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_2, B => \rc_shift[5]_net_1\, Y => 
        \rc_shift_30[4]_net_1\);
    
    \sd_ctl_p.sa_5[2]\ : CFG4
      generic map(INIT => x"C840")

      port map(A => act, B => sa_5_sn_N_4_mux, C => raddr(2), D
         => raddr(12), Y => sa_5_2);
    
    \pcable_shift_RNO[4]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[5]_net_1\, B => dorw(2), C => 
        bcount(2), Y => \pcable_shift_13[4]\);
    
    \rwable_shift[4]\ : SLE
      port map(D => \rwable_shift_7[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[4]_net_1\);
    
    \rc_shift_30[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_2, B => \rc_shift[2]_net_1\, Y => 
        \rc_shift_30[1]_net_1\);
    
    \actable_shift_57_m2[4]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[5]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[4]_net_1\);
    
    \sd_ctl_p.sa_5_1[1]\ : CFG3
      generic map(INIT => x"47")

      port map(A => raddr(11), B => act, C => raddr(1), Y => 
        \sa_5_1[1]\);
    
    \bterm_p.un4_bdzero_0_a2_RNI11LK\ : CFG4
      generic map(INIT => x"C084")

      port map(A => \CO1\, B => un4_bdzero, C => bdcnt(3), D => 
        bdcnt(2), Y => bdcnt_6_3);
    
    \actable_shift_57[12]\ : CFG4
      generic map(INIT => x"0FEE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[12]_net_1\, C => active(2), D => 
        refresh, Y => \actable_shift_57[12]_net_1\);
    
    \bterm_p.bdcnt_6_iv_0_m2[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => un14_rw, B => bdzero, C => rw, Y => N_68);
    
    \actable_shift[2]\ : SLE
      port map(D => \actable_shift_57[2]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[2]_net_1\);
    
    \actable_shift[7]\ : SLE
      port map(D => \actable_shift_57[7]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[7]_net_1\);
    
    CO1 : CFG2
      generic map(INIT => x"E")

      port map(A => bdcnt(0), B => bdcnt(1), Y => \CO1\);
    
    \act_p.3.un197_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => rwable_3, B => lnht_cmd(3), C => 
        un197_rdwr_cmd_0_a2_1, D => N_130, Y => \un197_rdwr_cmd\);
    
    \un1_mode_cmd\ : CFG3
      generic map(INIT => x"04")

      port map(A => prch_cmd, B => mode_cmd, C => rfsh_cmd, Y => 
        un1_mode_cmd);
    
    actable : SLE
      port map(D => actable_6, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => actable_2);
    
    un1_pch_3 : CFG4
      generic map(INIT => x"0100")

      port map(A => bterm, B => pch, C => rw, D => un36_rw_i_0_3, 
        Y => \un1_pch_3_i\);
    
    \act_p.3.un217_rdwr_cmd_0_a2_RNI89HJ\ : CFG3
      generic map(INIT => x"FE")

      port map(A => pch, B => \un217_rdwr_cmd\, C => bterm_cmd, Y
         => N_77);
    
    un1_rw_11 : CFG3
      generic map(INIT => x"01")

      port map(A => bcount(0), B => bcount(2), C => un28_rw, Y
         => \un1_rw_11_i\);
    
    \pcable_shift_RNO[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[4]_net_1\, B => dorw(2), C => 
        bcount(2), Y => N_752_i);
    
    actable_shift_57_ss0 : CFG3
      generic map(INIT => x"B8")

      port map(A => mode, B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_ss0\);
    
    \sd_ctl_p.sa_5[3]\ : CFG4
      generic map(INIT => x"C840")

      port map(A => act, B => sa_5_sn_N_4_mux, C => raddr(3), D
         => raddr(13), Y => sa_5_3);
    
    actable_6_iv : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \actable_1_sqmuxa_2\, B => un1_goactive_4_i, 
        C => \actable_shift[0]_net_1\, D => \rc_shift[0]_net_1\, 
        Y => actable_6);
    
    \act_p.1.un113_rdwr_cmd_0_a2_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => dorw(1), B => rdwr_cmd(1), Y => 
        un113_rdwr_cmd_0_a2_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity openbank_2 is

    port( bcount     : in    std_logic_vector(2 downto 0);
          raddr      : in    std_logic_vector(22 downto 10);
          line_i_3   : out   std_logic_vector(11 downto 0);
          prch_0     : in    std_logic;
          dorw_0     : in    std_logic;
          actable_0  : out   std_logic;
          rwable_0   : out   std_logic;
          pcable_0   : out   std_logic;
          chip_i_3_0 : out   std_logic;
          active_0   : out   std_logic;
          goact_0    : in    std_logic;
          refresh    : in    std_logic;
          mode       : in    std_logic;
          act        : in    std_logic;
          read_cmd   : in    std_logic;
          precharge  : in    std_logic;
          cke        : in    std_logic;
          clk        : in    std_logic;
          reset_n    : in    std_logic
        );

end openbank_2;

architecture DEF_ARCH of openbank_2 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \actable_shift[8]_net_1\, GND_net_1, 
        \actable_shift_57[8]_net_1\, VCC_net_1, 
        \actable_shift[9]_net_1\, \actable_shift_57[9]_net_1\, 
        \actable_shift[10]_net_1\, \actable_shift_57[10]_net_1\, 
        \actable_shift[11]_net_1\, \actable_shift_57[11]_net_1\, 
        \actable_shift[12]_net_1\, \actable_shift_57[12]_net_1\, 
        \pcable_shift[3]_net_1\, N_775_i, \pcable_shift[4]_net_1\, 
        \pcable_shift_13[4]\, \pcable_shift[5]_net_1\, 
        \pcable_shift_13[5]\, \pcable_shift[6]_net_1\, N_773_i, 
        \pcable_shift[7]_net_1\, \pcable_shift_13[7]\, 
        \pcable_shift[8]_net_1\, \pcable_shift_0_sqmuxa_i\, 
        \rc_shift[7]_net_1\, \rc_shift_30[7]_net_1\, 
        \rwable_shift[0]_net_1\, \rwable_shift_7[0]\, 
        \rwable_shift[1]_net_1\, \rwable_shift_7[1]\, 
        \rwable_shift[2]_net_1\, \rwable_shift_7[2]\, 
        \rwable_shift[3]_net_1\, \rwable_shift_7[3]\, 
        \rwable_shift[4]_net_1\, \rwable_shift_7[4]\, 
        \actable_shift[0]_net_1\, \actable_shift_57[0]_net_1\, 
        \actable_shift[1]_net_1\, \actable_shift_57[1]_net_1\, 
        \actable_shift[2]_net_1\, \actable_shift_57[2]_net_1\, 
        \actable_shift[3]_net_1\, \actable_shift_57[3]_net_1\, 
        \actable_shift[4]_net_1\, \actable_shift_57[4]_net_1\, 
        \actable_shift[5]_net_1\, \actable_shift_57[5]_net_1\, 
        \actable_shift[6]_net_1\, \actable_shift_57[6]_net_1\, 
        \actable_shift[7]_net_1\, \actable_shift_57[7]_net_1\, 
        \rc_shift[0]_net_1\, \rc_shift_30[0]_net_1\, 
        \rc_shift[1]_net_1\, \rc_shift_30[1]_net_1\, 
        \rc_shift[2]_net_1\, \rc_shift_30[2]_net_1\, 
        \rc_shift[3]_net_1\, \rc_shift_30[3]_net_1\, 
        \rc_shift[4]_net_1\, \rc_shift_30[4]_net_1\, 
        \rc_shift[5]_net_1\, \rc_shift_30[5]_net_1\, 
        \rc_shift[6]_net_1\, \rc_shift_30[6]_net_1\, \active_0\, 
        un36_dopch, \prev_cmd_read\, prev_cmd_read_1_2, N_774_i, 
        rwable_int_3, actable_6, un5_dopch_i, N_780, 
        \un1_goactive_4_1\, \actable_1_sqmuxa_2\, 
        un1_goactive_4_i, actable_shift_57_sm0, 
        \actable_shift_57_m2[12]_net_1\, \actable_shift_57_ss0\, 
        \actable_shift_57_m2[11]_net_1\, 
        \actable_shift_57_m2[10]_net_1\, 
        \actable_shift_57_m2[9]_net_1\, 
        \actable_shift_57_m2[8]_net_1\, 
        \actable_shift_57_m2[7]_net_1\, 
        \actable_shift_57_m2[6]_net_1\, 
        \actable_shift_57_m2[5]_net_1\, 
        \actable_shift_57_m2[4]_net_1\, 
        \actable_shift_57_m2[3]_net_1\, 
        \actable_shift_57_m2[2]_net_1\, 
        \actable_shift_57_m2[1]_net_1\ : std_logic;

begin 

    active_0 <= \active_0\;

    \rc_shift_30[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[5]_net_1\, Y => 
        \rc_shift_30[4]_net_1\);
    
    \rc_shift_30[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[4]_net_1\, Y => 
        \rc_shift_30[3]_net_1\);
    
    \actable_shift_57[1]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[1]_net_1\, Y => 
        \actable_shift_57[1]_net_1\);
    
    \pcable_shift[5]\ : SLE
      port map(D => \pcable_shift_13[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[5]_net_1\);
    
    \actable_shift_57[8]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[8]_net_1\, C => 
        \actable_shift[9]_net_1\, D => refresh, Y => 
        \actable_shift_57[8]_net_1\);
    
    \line[3]\ : SLE
      port map(D => raddr(13), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(3));
    
    \rc_shift[7]\ : SLE
      port map(D => \rc_shift_30[7]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[7]_net_1\);
    
    \pcable_shift[7]\ : SLE
      port map(D => \pcable_shift_13[7]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[7]_net_1\);
    
    \rc_shift_30[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[3]_net_1\, Y => 
        \rc_shift_30[2]_net_1\);
    
    \line[10]\ : SLE
      port map(D => raddr(20), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(10));
    
    \rc_shift_30[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => cke, Y => 
        \rc_shift_30[7]_net_1\);
    
    \actable_shift_57[4]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[4]_net_1\, Y => 
        \actable_shift_57[4]_net_1\);
    
    \rc_shift_30[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[1]_net_1\, Y => 
        \rc_shift_30[0]_net_1\);
    
    \rc_shift[3]\ : SLE
      port map(D => \rc_shift_30[3]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[3]_net_1\);
    
    \pcable_shift_RNO[7]\ : CFG4
      generic map(INIT => x"2AAA")

      port map(A => \pcable_shift[8]_net_1\, B => dorw_0, C => 
        bcount(1), D => bcount(2), Y => \pcable_shift_13[7]\);
    
    \actable_shift_57[0]\ : CFG4
      generic map(INIT => x"00EA")

      port map(A => un5_dopch_i, B => \actable_shift_57_ss0\, C
         => \actable_shift[1]_net_1\, D => refresh, Y => 
        \actable_shift_57[0]_net_1\);
    
    \actable_shift[5]\ : SLE
      port map(D => \actable_shift_57[5]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[5]_net_1\);
    
    actable : SLE
      port map(D => actable_6, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => actable_0);
    
    \rc_shift[0]\ : SLE
      port map(D => \rc_shift_30[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[0]_net_1\);
    
    \pcable_shift_RNO[5]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[6]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[5]\);
    
    \actable_shift_57_m2[10]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[11]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[10]_net_1\);
    
    \actable_shift[8]\ : SLE
      port map(D => \actable_shift_57[8]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[8]_net_1\);
    
    \actable_shift[0]\ : SLE
      port map(D => \actable_shift_57[0]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[0]_net_1\);
    
    prev_cmd_read : SLE
      port map(D => prev_cmd_read_1_2, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \prev_cmd_read\);
    
    actable_shift_57_ss0 : CFG3
      generic map(INIT => x"B8")

      port map(A => mode, B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_ss0\);
    
    \rw_p.rwable_shift_7[4]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => \active_0\, B => goact_0, C => un5_dopch_i, Y
         => \rwable_shift_7[4]\);
    
    \actable_shift[10]\ : SLE
      port map(D => \actable_shift_57[10]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[10]_net_1\);
    
    prev_cmd_read_1 : CFG3
      generic map(INIT => x"D8")

      port map(A => dorw_0, B => read_cmd, C => \prev_cmd_read\, 
        Y => prev_cmd_read_1_2);
    
    \pcable_shift[4]\ : SLE
      port map(D => \pcable_shift_13[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[4]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \actable_shift[12]\ : SLE
      port map(D => \actable_shift_57[12]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[12]_net_1\);
    
    \actable_shift[7]\ : SLE
      port map(D => \actable_shift_57[7]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[7]_net_1\);
    
    rwable_int : SLE
      port map(D => rwable_int_3, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rwable_0);
    
    pcable_int : SLE
      port map(D => N_774_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => pcable_0);
    
    \rw_p.rwable_int_3_iv\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[0]_net_1\, Y => rwable_int_3);
    
    \actable_shift[9]\ : SLE
      port map(D => \actable_shift_57[9]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[9]_net_1\);
    
    \actable_shift_57_m2[8]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[9]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[8]_net_1\);
    
    \actable_shift_57[3]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[3]_net_1\, Y => 
        \actable_shift_57[3]_net_1\);
    
    \rwable_shift[2]\ : SLE
      port map(D => \rwable_shift_7[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[2]_net_1\);
    
    \actable_shift[3]\ : SLE
      port map(D => \actable_shift_57[3]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[3]_net_1\);
    
    \line[5]\ : SLE
      port map(D => raddr(15), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(5));
    
    \rc_shift[4]\ : SLE
      port map(D => \rc_shift_30[4]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[4]_net_1\);
    
    \rw_p.rwable_shift_7[1]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[2]_net_1\, Y => \rwable_shift_7[1]\);
    
    \rwable_shift[4]\ : SLE
      port map(D => \rwable_shift_7[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[4]_net_1\);
    
    \actable_shift_57_m2[7]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[8]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[7]_net_1\);
    
    \pcable_shift[3]\ : SLE
      port map(D => N_775_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[3]_net_1\);
    
    \actable_shift[4]\ : SLE
      port map(D => \actable_shift_57[4]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[4]_net_1\);
    
    \actable_shift[11]\ : SLE
      port map(D => \actable_shift_57[11]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[11]_net_1\);
    
    \actable_shift_57[7]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[7]_net_1\, C => 
        \actable_shift[8]_net_1\, D => refresh, Y => 
        \actable_shift_57[7]_net_1\);
    
    \actable_shift[1]\ : SLE
      port map(D => \actable_shift_57[1]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \pcable_shift_RNO[4]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[5]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[4]\);
    
    \actable_shift_57_m2[4]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[5]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[4]_net_1\);
    
    \actable_shift_57_m2[11]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[12]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[11]_net_1\);
    
    un5_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => precharge, B => prch_0, Y => un5_dopch_i);
    
    \line[2]\ : SLE
      port map(D => raddr(12), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(2));
    
    \chip[0]\ : SLE
      port map(D => raddr(22), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => chip_i_3_0);
    
    \pcable_shift_RNO[6]\ : CFG4
      generic map(INIT => x"02AA")

      port map(A => \pcable_shift[7]_net_1\, B => bcount(0), C
         => bcount(1), D => N_780, Y => N_773_i);
    
    \rc_shift[1]\ : SLE
      port map(D => \rc_shift_30[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[1]_net_1\);
    
    \rc_shift[6]\ : SLE
      port map(D => \rc_shift_30[6]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[6]_net_1\);
    
    \line[4]\ : SLE
      port map(D => raddr(14), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(4));
    
    \rw_p.rwable_shift_7[2]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[3]_net_1\, Y => \rwable_shift_7[2]\);
    
    \actable_shift_57[10]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[10]_net_1\, C => 
        \actable_shift[11]_net_1\, D => refresh, Y => 
        \actable_shift_57[10]_net_1\);
    
    \actable_shift_57_m2[6]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[7]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[6]_net_1\);
    
    actable_1_sqmuxa_2 : CFG4
      generic map(INIT => x"0008")

      port map(A => \rc_shift[0]_net_1\, B => mode, C => refresh, 
        D => un5_dopch_i, Y => \actable_1_sqmuxa_2\);
    
    \line[11]\ : SLE
      port map(D => raddr(21), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(11));
    
    pcable_int_RNO : CFG4
      generic map(INIT => x"0E04")

      port map(A => \prev_cmd_read\, B => \pcable_shift[3]_net_1\, 
        C => dorw_0, D => \pcable_shift[4]_net_1\, Y => N_774_i);
    
    \rc_shift_30[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[2]_net_1\, Y => 
        \rc_shift_30[1]_net_1\);
    
    \actable_shift_57_m2[12]\ : CFG3
      generic map(INIT => x"54")

      port map(A => \active_0\, B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_m2[12]_net_1\);
    
    \actable_shift_57_m2[3]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[4]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[3]_net_1\);
    
    \line[9]\ : SLE
      port map(D => raddr(19), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(9));
    
    \line[1]\ : SLE
      port map(D => raddr(11), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(1));
    
    \actable_shift_57[6]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[6]_net_1\, C => 
        \actable_shift[7]_net_1\, D => refresh, Y => 
        \actable_shift_57[6]_net_1\);
    
    \actable_shift_57_m2[1]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[2]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[1]_net_1\);
    
    \pcable_shift[8]\ : SLE
      port map(D => \pcable_shift_0_sqmuxa_i\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[8]_net_1\);
    
    \rw_p.rwable_shift_7[0]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[1]_net_1\, Y => \rwable_shift_7[0]\);
    
    \rc_shift[5]\ : SLE
      port map(D => \rc_shift_30[5]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[5]_net_1\);
    
    \rc_shift_30[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[6]_net_1\, Y => 
        \rc_shift_30[5]_net_1\);
    
    \pcable_shift[6]\ : SLE
      port map(D => N_773_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[6]_net_1\);
    
    un1_goactive_4_1 : CFG4
      generic map(INIT => x"0031")

      port map(A => act, B => goact_0, C => \active_0\, D => mode, 
        Y => \un1_goactive_4_1\);
    
    \line[8]\ : SLE
      port map(D => raddr(18), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(8));
    
    active_int : SLE
      port map(D => goact_0, CLK => clk, EN => un36_dopch, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \active_0\);
    
    \actable_shift_57_m2[9]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[10]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[9]_net_1\);
    
    \rw_p.rwable_shift_7[3]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[4]_net_1\, Y => \rwable_shift_7[3]\);
    
    \line[0]\ : SLE
      port map(D => raddr(10), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(0));
    
    \rwable_shift[1]\ : SLE
      port map(D => \rwable_shift_7[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[1]_net_1\);
    
    un1_pcable_shift_3_sqmuxa_i_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => bcount(2), B => dorw_0, Y => N_780);
    
    actable_6_iv : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \actable_1_sqmuxa_2\, B => un1_goactive_4_i, 
        C => \actable_shift[0]_net_1\, D => \rc_shift[0]_net_1\, 
        Y => actable_6);
    
    \rc_shift[2]\ : SLE
      port map(D => \rc_shift_30[2]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[2]_net_1\);
    
    \line[7]\ : SLE
      port map(D => raddr(17), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(7));
    
    \actable_shift_57[9]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[9]_net_1\, C => 
        \actable_shift[10]_net_1\, D => refresh, Y => 
        \actable_shift_57[9]_net_1\);
    
    \actable_shift_57[11]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[11]_net_1\, C => 
        \actable_shift[12]_net_1\, D => refresh, Y => 
        \actable_shift_57[11]_net_1\);
    
    \rc_shift_30[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[7]_net_1\, Y => 
        \rc_shift_30[6]_net_1\);
    
    \actable_shift_57[2]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[2]_net_1\, Y => 
        \actable_shift_57[2]_net_1\);
    
    \actable_shift_57[12]\ : CFG4
      generic map(INIT => x"0FEE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[12]_net_1\, C => \active_0\, D => 
        refresh, Y => \actable_shift_57[12]_net_1\);
    
    \actable_shift[6]\ : SLE
      port map(D => \actable_shift_57[6]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[6]_net_1\);
    
    un7_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => un5_dopch_i, B => goact_0, Y => un36_dopch);
    
    \pcable_shift_RNO[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[4]_net_1\, B => dorw_0, C => 
        bcount(2), Y => N_775_i);
    
    un1_goactive_4 : CFG3
      generic map(INIT => x"10")

      port map(A => refresh, B => un5_dopch_i, C => 
        \un1_goactive_4_1\, Y => un1_goactive_4_i);
    
    actable_shift_57_m2s2 : CFG4
      generic map(INIT => x"FF02")

      port map(A => act, B => goact_0, C => \active_0\, D => mode, 
        Y => actable_shift_57_sm0);
    
    \rwable_shift[0]\ : SLE
      port map(D => \rwable_shift_7[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[0]_net_1\);
    
    \actable_shift_57_m2[2]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[3]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[2]_net_1\);
    
    \rwable_shift[3]\ : SLE
      port map(D => \rwable_shift_7[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[3]_net_1\);
    
    pcable_shift_0_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bcount(1), B => bcount(2), C => dorw_0, D => 
        bcount(0), Y => \pcable_shift_0_sqmuxa_i\);
    
    \actable_shift_57_m2[5]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[6]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[5]_net_1\);
    
    \actable_shift[2]\ : SLE
      port map(D => \actable_shift_57[2]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[2]_net_1\);
    
    \actable_shift_57[5]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[5]_net_1\, Y => 
        \actable_shift_57[5]_net_1\);
    
    \line[6]\ : SLE
      port map(D => raddr(16), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_3(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity openbank_0 is

    port( bcount              : in    std_logic_vector(2 downto 0);
          raddr               : in    std_logic_vector(22 downto 10);
          line_i_1            : out   std_logic_vector(11 downto 0);
          sa_5_0              : out   std_logic;
          sa_5_2              : out   std_logic;
          prch_0              : in    std_logic;
          dorw_0              : in    std_logic;
          actable_0           : out   std_logic;
          rwable_0            : out   std_logic;
          pcable_0            : out   std_logic;
          chip_i_1_0          : out   std_logic;
          active_0            : out   std_logic;
          goact_0             : in    std_logic;
          pch                 : in    std_logic;
          un8_precharge       : in    std_logic;
          act                 : in    std_logic;
          read_cmd            : in    std_logic;
          precharge           : in    std_logic;
          cas_n_1             : out   std_logic;
          un1_precharge_5_i_0 : in    std_logic;
          ras_n_1             : out   std_logic;
          un1_precharge_3_i_0 : in    std_logic;
          cke                 : in    std_logic;
          mode                : in    std_logic;
          refresh             : in    std_logic;
          clk                 : in    std_logic;
          reset_n             : in    std_logic
        );

end openbank_0;

architecture DEF_ARCH of openbank_0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \actable_shift[8]_net_1\, GND_net_1, 
        \actable_shift_57[8]_net_1\, VCC_net_1, 
        \actable_shift[9]_net_1\, \actable_shift_57[9]_net_1\, 
        \actable_shift[10]_net_1\, \actable_shift_57[10]_net_1\, 
        \actable_shift[11]_net_1\, \actable_shift_57[11]_net_1\, 
        \actable_shift[12]_net_1\, \actable_shift_57[12]_net_1\, 
        \pcable_shift[3]_net_1\, N_759_i, \pcable_shift[4]_net_1\, 
        \pcable_shift_13[4]\, \pcable_shift[5]_net_1\, 
        \pcable_shift_13[5]\, \pcable_shift[6]_net_1\, N_757_i, 
        \pcable_shift[7]_net_1\, \pcable_shift_13[7]\, 
        \pcable_shift[8]_net_1\, \pcable_shift_0_sqmuxa_i\, 
        \rc_shift[7]_net_1\, \rc_shift_30[7]_net_1\, 
        \rwable_shift[0]_net_1\, \rwable_shift_7[0]\, 
        \rwable_shift[1]_net_1\, \rwable_shift_7[1]\, 
        \rwable_shift[2]_net_1\, \rwable_shift_7[2]\, 
        \rwable_shift[3]_net_1\, \rwable_shift_7[3]\, 
        \rwable_shift[4]_net_1\, \rwable_shift_7[4]\, 
        \actable_shift[0]_net_1\, \actable_shift_57[0]_net_1\, 
        \actable_shift[1]_net_1\, \actable_shift_57[1]_net_1\, 
        \actable_shift[2]_net_1\, \actable_shift_57[2]_net_1\, 
        \actable_shift[3]_net_1\, \actable_shift_57[3]_net_1\, 
        \actable_shift[4]_net_1\, \actable_shift_57[4]_net_1\, 
        \actable_shift[5]_net_1\, \actable_shift_57[5]_net_1\, 
        \actable_shift[6]_net_1\, \actable_shift_57[6]_net_1\, 
        \actable_shift[7]_net_1\, \actable_shift_57[7]_net_1\, 
        \rc_shift[0]_net_1\, \rc_shift_30[0]_net_1\, 
        \rc_shift[1]_net_1\, \rc_shift_30[1]_net_1\, 
        \rc_shift[2]_net_1\, \rc_shift_30[2]_net_1\, 
        \rc_shift[3]_net_1\, \rc_shift_30[3]_net_1\, 
        \rc_shift[4]_net_1\, \rc_shift_30[4]_net_1\, 
        \rc_shift[5]_net_1\, \rc_shift_30[5]_net_1\, 
        \rc_shift[6]_net_1\, \rc_shift_30[6]_net_1\, \active_0\, 
        un36_dopch, \prev_cmd_read\, prev_cmd_read_1_0, N_758_i, 
        rwable_int_3, actable_6, un5_dopch_i, 
        \actable_1_sqmuxa_2\, N_764, \un1_goactive_4_1\, 
        \un2_domode\, un1_goactive_4_i, \actable_shift_5_sqmuxa\, 
        \actable_shift_57_m2[11]_net_1\, 
        \actable_shift_57_m2[10]_net_1\, 
        \actable_shift_57_m2[9]_net_1\, 
        \actable_shift_57_m2[8]_net_1\, 
        \actable_shift_57_m2[7]_net_1\, 
        \actable_shift_57_m2[6]_net_1\, 
        \actable_shift_57_m2[5]_net_1\, 
        \actable_shift_57_m2[4]_net_1\, 
        \actable_shift_57_m2[3]_net_1\, 
        \actable_shift_57_m2[2]_net_1\, 
        \actable_shift_57_m2[1]_net_1\, \actable_shift_57_ss0\, 
        \actable_shift_57_m2[12]_net_1\ : std_logic;

begin 

    active_0 <= \active_0\;

    \rc_shift_30[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[5]_net_1\, Y => 
        \rc_shift_30[4]_net_1\);
    
    \rc_shift_30[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[4]_net_1\, Y => 
        \rc_shift_30[3]_net_1\);
    
    \actable_shift_57[1]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[1]_net_1\, Y => 
        \actable_shift_57[1]_net_1\);
    
    \pcable_shift[5]\ : SLE
      port map(D => \pcable_shift_13[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[5]_net_1\);
    
    \actable_shift_57[8]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[8]_net_1\, C => 
        \actable_shift[9]_net_1\, D => refresh, Y => 
        \actable_shift_57[8]_net_1\);
    
    \line[3]\ : SLE
      port map(D => raddr(13), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(3));
    
    \rc_shift[7]\ : SLE
      port map(D => \rc_shift_30[7]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[7]_net_1\);
    
    \pcable_shift[7]\ : SLE
      port map(D => \pcable_shift_13[7]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[7]_net_1\);
    
    \rc_shift_30[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[3]_net_1\, Y => 
        \rc_shift_30[2]_net_1\);
    
    \line[10]\ : SLE
      port map(D => raddr(20), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(10));
    
    \rc_shift_30[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => cke, Y => 
        \rc_shift_30[7]_net_1\);
    
    \actable_shift_57[4]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[4]_net_1\, Y => 
        \actable_shift_57[4]_net_1\);
    
    \sd_ctl_p.sa_5[9]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => act, B => un8_precharge, C => pch, D => 
        raddr(19), Y => sa_5_0);
    
    \rc_shift_30[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[1]_net_1\, Y => 
        \rc_shift_30[0]_net_1\);
    
    \rc_shift[3]\ : SLE
      port map(D => \rc_shift_30[3]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[3]_net_1\);
    
    \pcable_shift_RNO[7]\ : CFG4
      generic map(INIT => x"2AAA")

      port map(A => \pcable_shift[8]_net_1\, B => dorw_0, C => 
        bcount(1), D => bcount(2), Y => \pcable_shift_13[7]\);
    
    \actable_shift_57[0]\ : CFG4
      generic map(INIT => x"00EA")

      port map(A => un5_dopch_i, B => \actable_shift_57_ss0\, C
         => \actable_shift[1]_net_1\, D => refresh, Y => 
        \actable_shift_57[0]_net_1\);
    
    \actable_shift[5]\ : SLE
      port map(D => \actable_shift_57[5]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[5]_net_1\);
    
    actable : SLE
      port map(D => actable_6, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => actable_0);
    
    \rc_shift[0]\ : SLE
      port map(D => \rc_shift_30[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[0]_net_1\);
    
    \pcable_shift_RNO[5]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[6]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[5]\);
    
    \actable_shift_57_m2[10]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[11]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[10]_net_1\);
    
    \actable_shift[8]\ : SLE
      port map(D => \actable_shift_57[8]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[8]_net_1\);
    
    \actable_shift[0]\ : SLE
      port map(D => \actable_shift_57[0]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[0]_net_1\);
    
    prev_cmd_read : SLE
      port map(D => prev_cmd_read_1_0, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \prev_cmd_read\);
    
    actable_shift_57_ss0 : CFG4
      generic map(INIT => x"F0E4")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => mode, D => \un2_domode\, Y => 
        \actable_shift_57_ss0\);
    
    \rw_p.rwable_shift_7[4]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => \active_0\, B => goact_0, C => un5_dopch_i, Y
         => \rwable_shift_7[4]\);
    
    \actable_shift[10]\ : SLE
      port map(D => \actable_shift_57[10]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[10]_net_1\);
    
    prev_cmd_read_1 : CFG3
      generic map(INIT => x"D8")

      port map(A => dorw_0, B => read_cmd, C => \prev_cmd_read\, 
        Y => prev_cmd_read_1_0);
    
    \pcable_shift[4]\ : SLE
      port map(D => \pcable_shift_13[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[4]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \actable_shift[12]\ : SLE
      port map(D => \actable_shift_57[12]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[12]_net_1\);
    
    \sd_ctl_p.sa_5[11]\ : CFG4
      generic map(INIT => x"0200")

      port map(A => act, B => un8_precharge, C => pch, D => 
        raddr(21), Y => sa_5_2);
    
    \actable_shift[7]\ : SLE
      port map(D => \actable_shift_57[7]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[7]_net_1\);
    
    rwable_int : SLE
      port map(D => rwable_int_3, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rwable_0);
    
    pcable_int : SLE
      port map(D => N_758_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => pcable_0);
    
    un2_domode : CFG3
      generic map(INIT => x"04")

      port map(A => un5_dopch_i, B => mode, C => refresh, Y => 
        \un2_domode\);
    
    \rw_p.rwable_int_3_iv\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[0]_net_1\, Y => rwable_int_3);
    
    \actable_shift[9]\ : SLE
      port map(D => \actable_shift_57[9]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[9]_net_1\);
    
    \actable_shift_57_m2[8]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[9]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[8]_net_1\);
    
    \actable_shift_57[3]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[3]_net_1\, Y => 
        \actable_shift_57[3]_net_1\);
    
    \rwable_shift[2]\ : SLE
      port map(D => \rwable_shift_7[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[2]_net_1\);
    
    \actable_shift[3]\ : SLE
      port map(D => \actable_shift_57[3]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[3]_net_1\);
    
    \line[5]\ : SLE
      port map(D => raddr(15), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(5));
    
    actable_shift_5_sqmuxa : CFG4
      generic map(INIT => x"0002")

      port map(A => act, B => \active_0\, C => un5_dopch_i, D => 
        goact_0, Y => \actable_shift_5_sqmuxa\);
    
    \rc_shift[4]\ : SLE
      port map(D => \rc_shift_30[4]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[4]_net_1\);
    
    \rw_p.rwable_shift_7[1]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[2]_net_1\, Y => \rwable_shift_7[1]\);
    
    \rwable_shift[4]\ : SLE
      port map(D => \rwable_shift_7[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[4]_net_1\);
    
    \actable_shift_57_m2[7]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[8]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[7]_net_1\);
    
    \pcable_shift[3]\ : SLE
      port map(D => N_759_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[3]_net_1\);
    
    \actable_shift[4]\ : SLE
      port map(D => \actable_shift_57[4]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[4]_net_1\);
    
    \actable_shift[11]\ : SLE
      port map(D => \actable_shift_57[11]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[11]_net_1\);
    
    \actable_shift_57[7]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[7]_net_1\, C => 
        \actable_shift[8]_net_1\, D => refresh, Y => 
        \actable_shift_57[7]_net_1\);
    
    \actable_shift[1]\ : SLE
      port map(D => \actable_shift_57[1]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sd_ctl_p.cas_n_1_0_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => un1_precharge_5_i_0, B => refresh, Y => 
        cas_n_1);
    
    \pcable_shift_RNO[4]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[5]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[4]\);
    
    \actable_shift_57_m2[4]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[5]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[4]_net_1\);
    
    \actable_shift_57_m2[11]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[12]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[11]_net_1\);
    
    un5_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => precharge, B => prch_0, Y => un5_dopch_i);
    
    \line[2]\ : SLE
      port map(D => raddr(12), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(2));
    
    \chip[0]\ : SLE
      port map(D => raddr(22), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => chip_i_1_0);
    
    \pcable_shift_RNO[6]\ : CFG4
      generic map(INIT => x"02AA")

      port map(A => \pcable_shift[7]_net_1\, B => bcount(0), C
         => bcount(1), D => N_764, Y => N_757_i);
    
    \rc_shift[1]\ : SLE
      port map(D => \rc_shift_30[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[1]_net_1\);
    
    \rc_shift[6]\ : SLE
      port map(D => \rc_shift_30[6]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[6]_net_1\);
    
    \line[4]\ : SLE
      port map(D => raddr(14), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(4));
    
    \rw_p.rwable_shift_7[2]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[3]_net_1\, Y => \rwable_shift_7[2]\);
    
    \actable_shift_57[10]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[10]_net_1\, C => 
        \actable_shift[11]_net_1\, D => refresh, Y => 
        \actable_shift_57[10]_net_1\);
    
    \actable_shift_57_m2[6]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[7]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[6]_net_1\);
    
    actable_1_sqmuxa_2 : CFG4
      generic map(INIT => x"1000")

      port map(A => refresh, B => un5_dopch_i, C => 
        \rc_shift[0]_net_1\, D => mode, Y => \actable_1_sqmuxa_2\);
    
    \line[11]\ : SLE
      port map(D => raddr(21), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(11));
    
    pcable_int_RNO : CFG4
      generic map(INIT => x"0E04")

      port map(A => \prev_cmd_read\, B => \pcable_shift[3]_net_1\, 
        C => dorw_0, D => \pcable_shift[4]_net_1\, Y => N_758_i);
    
    \rc_shift_30[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[2]_net_1\, Y => 
        \rc_shift_30[1]_net_1\);
    
    \actable_shift_57_m2[12]\ : CFG4
      generic map(INIT => x"0F0E")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \active_0\, D => \un2_domode\, Y
         => \actable_shift_57_m2[12]_net_1\);
    
    \actable_shift_57_m2[3]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[4]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[3]_net_1\);
    
    \line[9]\ : SLE
      port map(D => raddr(19), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(9));
    
    \line[1]\ : SLE
      port map(D => raddr(11), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(1));
    
    \actable_shift_57[6]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[6]_net_1\, C => 
        \actable_shift[7]_net_1\, D => refresh, Y => 
        \actable_shift_57[6]_net_1\);
    
    \actable_shift_57_m2[1]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[2]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[1]_net_1\);
    
    \pcable_shift[8]\ : SLE
      port map(D => \pcable_shift_0_sqmuxa_i\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[8]_net_1\);
    
    \rw_p.rwable_shift_7[0]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[1]_net_1\, Y => \rwable_shift_7[0]\);
    
    \rc_shift[5]\ : SLE
      port map(D => \rc_shift_30[5]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[5]_net_1\);
    
    \rc_shift_30[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[6]_net_1\, Y => 
        \rc_shift_30[5]_net_1\);
    
    \sd_ctl_p.ras_n_1_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_precharge_3_i_0, B => refresh, Y => 
        ras_n_1);
    
    \pcable_shift[6]\ : SLE
      port map(D => N_757_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[6]_net_1\);
    
    un1_goactive_4_1 : CFG4
      generic map(INIT => x"0031")

      port map(A => act, B => goact_0, C => \active_0\, D => mode, 
        Y => \un1_goactive_4_1\);
    
    \line[8]\ : SLE
      port map(D => raddr(18), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(8));
    
    active_int : SLE
      port map(D => goact_0, CLK => clk, EN => un36_dopch, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \active_0\);
    
    \actable_shift_57_m2[9]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[10]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[9]_net_1\);
    
    \rw_p.rwable_shift_7[3]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[4]_net_1\, Y => \rwable_shift_7[3]\);
    
    \line[0]\ : SLE
      port map(D => raddr(10), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(0));
    
    \rwable_shift[1]\ : SLE
      port map(D => \rwable_shift_7[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[1]_net_1\);
    
    un1_pcable_shift_3_sqmuxa_i_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => bcount(2), B => dorw_0, Y => N_764);
    
    actable_6_iv : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \actable_1_sqmuxa_2\, B => un1_goactive_4_i, 
        C => \actable_shift[0]_net_1\, D => \rc_shift[0]_net_1\, 
        Y => actable_6);
    
    \rc_shift[2]\ : SLE
      port map(D => \rc_shift_30[2]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[2]_net_1\);
    
    \line[7]\ : SLE
      port map(D => raddr(17), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(7));
    
    \actable_shift_57[9]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[9]_net_1\, C => 
        \actable_shift[10]_net_1\, D => refresh, Y => 
        \actable_shift_57[9]_net_1\);
    
    \actable_shift_57[11]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[11]_net_1\, C => 
        \actable_shift[12]_net_1\, D => refresh, Y => 
        \actable_shift_57[11]_net_1\);
    
    \rc_shift_30[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[7]_net_1\, Y => 
        \rc_shift_30[6]_net_1\);
    
    \actable_shift_57[2]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[2]_net_1\, Y => 
        \actable_shift_57[2]_net_1\);
    
    \actable_shift_57[12]\ : CFG4
      generic map(INIT => x"0FEE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[12]_net_1\, C => \active_0\, D => 
        refresh, Y => \actable_shift_57[12]_net_1\);
    
    \actable_shift[6]\ : SLE
      port map(D => \actable_shift_57[6]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[6]_net_1\);
    
    un7_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => un5_dopch_i, B => goact_0, Y => un36_dopch);
    
    \pcable_shift_RNO[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[4]_net_1\, B => dorw_0, C => 
        bcount(2), Y => N_759_i);
    
    un1_goactive_4 : CFG3
      generic map(INIT => x"10")

      port map(A => refresh, B => un5_dopch_i, C => 
        \un1_goactive_4_1\, Y => un1_goactive_4_i);
    
    \rwable_shift[0]\ : SLE
      port map(D => \rwable_shift_7[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[0]_net_1\);
    
    \actable_shift_57_m2[2]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[3]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[2]_net_1\);
    
    \rwable_shift[3]\ : SLE
      port map(D => \rwable_shift_7[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[3]_net_1\);
    
    pcable_shift_0_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bcount(1), B => bcount(2), C => dorw_0, D => 
        bcount(0), Y => \pcable_shift_0_sqmuxa_i\);
    
    \actable_shift_57_m2[5]\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => \actable_shift_5_sqmuxa\, B => 
        un1_goactive_4_i, C => \actable_shift[6]_net_1\, D => 
        \un2_domode\, Y => \actable_shift_57_m2[5]_net_1\);
    
    \actable_shift[2]\ : SLE
      port map(D => \actable_shift_57[2]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[2]_net_1\);
    
    \actable_shift_57[5]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[5]_net_1\, Y => 
        \actable_shift_57[5]_net_1\);
    
    \line[6]\ : SLE
      port map(D => raddr(16), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_1(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity openbank_1 is

    port( bcount     : in    std_logic_vector(2 downto 0);
          raddr      : in    std_logic_vector(22 downto 10);
          line_i_0   : out   std_logic_vector(11 downto 0);
          prch_0     : in    std_logic;
          dorw_0     : in    std_logic;
          actable_0  : out   std_logic;
          rwable_0   : out   std_logic;
          pcable_0   : out   std_logic;
          chip_i_0_0 : out   std_logic;
          active_0   : out   std_logic;
          goact_0    : in    std_logic;
          refresh    : in    std_logic;
          mode       : in    std_logic;
          act        : in    std_logic;
          read_cmd   : in    std_logic;
          precharge  : in    std_logic;
          cke        : in    std_logic;
          clk        : in    std_logic;
          reset_n    : in    std_logic
        );

end openbank_1;

architecture DEF_ARCH of openbank_1 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \actable_shift[8]_net_1\, GND_net_1, 
        \actable_shift_57[8]_net_1\, VCC_net_1, 
        \actable_shift[9]_net_1\, \actable_shift_57[9]_net_1\, 
        \actable_shift[10]_net_1\, \actable_shift_57[10]_net_1\, 
        \actable_shift[11]_net_1\, \actable_shift_57[11]_net_1\, 
        \actable_shift[12]_net_1\, \actable_shift_57[12]_net_1\, 
        \pcable_shift[3]_net_1\, N_767_i, \pcable_shift[4]_net_1\, 
        \pcable_shift_13[4]\, \pcable_shift[5]_net_1\, 
        \pcable_shift_13[5]\, \pcable_shift[6]_net_1\, N_765_i, 
        \pcable_shift[7]_net_1\, \pcable_shift_13[7]\, 
        \pcable_shift[8]_net_1\, \pcable_shift_0_sqmuxa_i\, 
        \rc_shift[7]_net_1\, \rc_shift_30[7]_net_1\, 
        \rwable_shift[0]_net_1\, \rwable_shift_7[0]\, 
        \rwable_shift[1]_net_1\, \rwable_shift_7[1]\, 
        \rwable_shift[2]_net_1\, \rwable_shift_7[2]\, 
        \rwable_shift[3]_net_1\, \rwable_shift_7[3]\, 
        \rwable_shift[4]_net_1\, \rwable_shift_7[4]\, 
        \actable_shift[0]_net_1\, \actable_shift_57[0]_net_1\, 
        \actable_shift[1]_net_1\, \actable_shift_57[1]_net_1\, 
        \actable_shift[2]_net_1\, \actable_shift_57[2]_net_1\, 
        \actable_shift[3]_net_1\, \actable_shift_57[3]_net_1\, 
        \actable_shift[4]_net_1\, \actable_shift_57[4]_net_1\, 
        \actable_shift[5]_net_1\, \actable_shift_57[5]_net_1\, 
        \actable_shift[6]_net_1\, \actable_shift_57[6]_net_1\, 
        \actable_shift[7]_net_1\, \actable_shift_57[7]_net_1\, 
        \rc_shift[0]_net_1\, \rc_shift_30[0]_net_1\, 
        \rc_shift[1]_net_1\, \rc_shift_30[1]_net_1\, 
        \rc_shift[2]_net_1\, \rc_shift_30[2]_net_1\, 
        \rc_shift[3]_net_1\, \rc_shift_30[3]_net_1\, 
        \rc_shift[4]_net_1\, \rc_shift_30[4]_net_1\, 
        \rc_shift[5]_net_1\, \rc_shift_30[5]_net_1\, 
        \rc_shift[6]_net_1\, \rc_shift_30[6]_net_1\, \active_0\, 
        un36_dopch, \prev_cmd_read\, prev_cmd_read_1_1, N_766_i, 
        rwable_int_3, actable_6, un5_dopch_i, N_772, 
        \un1_goactive_4_1\, \actable_1_sqmuxa_2\, 
        un1_goactive_4_i, actable_shift_57_sm0, 
        \actable_shift_57_ss0\, \actable_shift_57_m2[1]_net_1\, 
        \actable_shift_57_m2[2]_net_1\, 
        \actable_shift_57_m2[3]_net_1\, 
        \actable_shift_57_m2[4]_net_1\, 
        \actable_shift_57_m2[5]_net_1\, 
        \actable_shift_57_m2[6]_net_1\, 
        \actable_shift_57_m2[7]_net_1\, 
        \actable_shift_57_m2[8]_net_1\, 
        \actable_shift_57_m2[9]_net_1\, 
        \actable_shift_57_m2[10]_net_1\, 
        \actable_shift_57_m2[11]_net_1\, 
        \actable_shift_57_m2[12]_net_1\ : std_logic;

begin 

    active_0 <= \active_0\;

    \rc_shift_30[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[5]_net_1\, Y => 
        \rc_shift_30[4]_net_1\);
    
    \rc_shift_30[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[4]_net_1\, Y => 
        \rc_shift_30[3]_net_1\);
    
    \actable_shift_57[1]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[1]_net_1\, Y => 
        \actable_shift_57[1]_net_1\);
    
    \pcable_shift[5]\ : SLE
      port map(D => \pcable_shift_13[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[5]_net_1\);
    
    \actable_shift_57[8]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[8]_net_1\, C => 
        \actable_shift[9]_net_1\, D => refresh, Y => 
        \actable_shift_57[8]_net_1\);
    
    \line[3]\ : SLE
      port map(D => raddr(13), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(3));
    
    \rc_shift[7]\ : SLE
      port map(D => \rc_shift_30[7]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[7]_net_1\);
    
    \pcable_shift[7]\ : SLE
      port map(D => \pcable_shift_13[7]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[7]_net_1\);
    
    \rc_shift_30[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[3]_net_1\, Y => 
        \rc_shift_30[2]_net_1\);
    
    \line[10]\ : SLE
      port map(D => raddr(20), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(10));
    
    \rc_shift_30[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => cke, Y => 
        \rc_shift_30[7]_net_1\);
    
    \actable_shift_57[4]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[4]_net_1\, Y => 
        \actable_shift_57[4]_net_1\);
    
    \rc_shift_30[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[1]_net_1\, Y => 
        \rc_shift_30[0]_net_1\);
    
    \rc_shift[3]\ : SLE
      port map(D => \rc_shift_30[3]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[3]_net_1\);
    
    \pcable_shift_RNO[7]\ : CFG4
      generic map(INIT => x"2AAA")

      port map(A => \pcable_shift[8]_net_1\, B => dorw_0, C => 
        bcount(1), D => bcount(2), Y => \pcable_shift_13[7]\);
    
    \actable_shift_57[0]\ : CFG4
      generic map(INIT => x"00EA")

      port map(A => un5_dopch_i, B => \actable_shift_57_ss0\, C
         => \actable_shift[1]_net_1\, D => refresh, Y => 
        \actable_shift_57[0]_net_1\);
    
    \actable_shift[5]\ : SLE
      port map(D => \actable_shift_57[5]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[5]_net_1\);
    
    actable : SLE
      port map(D => actable_6, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => actable_0);
    
    \rc_shift[0]\ : SLE
      port map(D => \rc_shift_30[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[0]_net_1\);
    
    \pcable_shift_RNO[5]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[6]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[5]\);
    
    \actable_shift_57_m2[10]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[11]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[10]_net_1\);
    
    \actable_shift[8]\ : SLE
      port map(D => \actable_shift_57[8]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[8]_net_1\);
    
    \actable_shift[0]\ : SLE
      port map(D => \actable_shift_57[0]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[0]_net_1\);
    
    prev_cmd_read : SLE
      port map(D => prev_cmd_read_1_1, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \prev_cmd_read\);
    
    actable_shift_57_ss0 : CFG3
      generic map(INIT => x"B8")

      port map(A => mode, B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_ss0\);
    
    \rw_p.rwable_shift_7[4]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => \active_0\, B => goact_0, C => un5_dopch_i, Y
         => \rwable_shift_7[4]\);
    
    \actable_shift[10]\ : SLE
      port map(D => \actable_shift_57[10]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[10]_net_1\);
    
    prev_cmd_read_1 : CFG3
      generic map(INIT => x"D8")

      port map(A => dorw_0, B => read_cmd, C => \prev_cmd_read\, 
        Y => prev_cmd_read_1_1);
    
    \pcable_shift[4]\ : SLE
      port map(D => \pcable_shift_13[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[4]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \actable_shift[12]\ : SLE
      port map(D => \actable_shift_57[12]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[12]_net_1\);
    
    \actable_shift[7]\ : SLE
      port map(D => \actable_shift_57[7]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[7]_net_1\);
    
    rwable_int : SLE
      port map(D => rwable_int_3, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rwable_0);
    
    pcable_int : SLE
      port map(D => N_766_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => pcable_0);
    
    \rw_p.rwable_int_3_iv\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[0]_net_1\, Y => rwable_int_3);
    
    \actable_shift[9]\ : SLE
      port map(D => \actable_shift_57[9]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[9]_net_1\);
    
    \actable_shift_57_m2[8]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[9]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[8]_net_1\);
    
    \actable_shift_57[3]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[3]_net_1\, Y => 
        \actable_shift_57[3]_net_1\);
    
    \rwable_shift[2]\ : SLE
      port map(D => \rwable_shift_7[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[2]_net_1\);
    
    \actable_shift[3]\ : SLE
      port map(D => \actable_shift_57[3]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[3]_net_1\);
    
    \line[5]\ : SLE
      port map(D => raddr(15), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(5));
    
    \rc_shift[4]\ : SLE
      port map(D => \rc_shift_30[4]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[4]_net_1\);
    
    \rw_p.rwable_shift_7[1]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[2]_net_1\, Y => \rwable_shift_7[1]\);
    
    \rwable_shift[4]\ : SLE
      port map(D => \rwable_shift_7[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[4]_net_1\);
    
    \actable_shift_57_m2[7]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[8]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[7]_net_1\);
    
    \pcable_shift[3]\ : SLE
      port map(D => N_767_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[3]_net_1\);
    
    \actable_shift[4]\ : SLE
      port map(D => \actable_shift_57[4]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[4]_net_1\);
    
    \actable_shift[11]\ : SLE
      port map(D => \actable_shift_57[11]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[11]_net_1\);
    
    \actable_shift_57[7]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[7]_net_1\, C => 
        \actable_shift[8]_net_1\, D => refresh, Y => 
        \actable_shift_57[7]_net_1\);
    
    \actable_shift[1]\ : SLE
      port map(D => \actable_shift_57[1]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \pcable_shift_RNO[4]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[5]_net_1\, B => dorw_0, C => 
        bcount(2), Y => \pcable_shift_13[4]\);
    
    \actable_shift_57_m2[4]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[5]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[4]_net_1\);
    
    \actable_shift_57_m2[11]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[12]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[11]_net_1\);
    
    un5_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => precharge, B => prch_0, Y => un5_dopch_i);
    
    \line[2]\ : SLE
      port map(D => raddr(12), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(2));
    
    \chip[0]\ : SLE
      port map(D => raddr(22), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => chip_i_0_0);
    
    \pcable_shift_RNO[6]\ : CFG4
      generic map(INIT => x"02AA")

      port map(A => \pcable_shift[7]_net_1\, B => bcount(0), C
         => bcount(1), D => N_772, Y => N_765_i);
    
    \rc_shift[1]\ : SLE
      port map(D => \rc_shift_30[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[1]_net_1\);
    
    \rc_shift[6]\ : SLE
      port map(D => \rc_shift_30[6]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[6]_net_1\);
    
    \line[4]\ : SLE
      port map(D => raddr(14), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(4));
    
    \rw_p.rwable_shift_7[2]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[3]_net_1\, Y => \rwable_shift_7[2]\);
    
    \actable_shift_57[10]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[10]_net_1\, C => 
        \actable_shift[11]_net_1\, D => refresh, Y => 
        \actable_shift_57[10]_net_1\);
    
    \actable_shift_57_m2[6]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[7]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[6]_net_1\);
    
    actable_1_sqmuxa_2 : CFG4
      generic map(INIT => x"0008")

      port map(A => \rc_shift[0]_net_1\, B => mode, C => refresh, 
        D => un5_dopch_i, Y => \actable_1_sqmuxa_2\);
    
    \line[11]\ : SLE
      port map(D => raddr(21), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(11));
    
    pcable_int_RNO : CFG4
      generic map(INIT => x"0E04")

      port map(A => \prev_cmd_read\, B => \pcable_shift[3]_net_1\, 
        C => dorw_0, D => \pcable_shift[4]_net_1\, Y => N_766_i);
    
    \rc_shift_30[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => goact_0, B => \rc_shift[2]_net_1\, Y => 
        \rc_shift_30[1]_net_1\);
    
    \actable_shift_57_m2[12]\ : CFG3
      generic map(INIT => x"54")

      port map(A => \active_0\, B => actable_shift_57_sm0, C => 
        un1_goactive_4_i, Y => \actable_shift_57_m2[12]_net_1\);
    
    \actable_shift_57_m2[3]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[4]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[3]_net_1\);
    
    \line[9]\ : SLE
      port map(D => raddr(19), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(9));
    
    \line[1]\ : SLE
      port map(D => raddr(11), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(1));
    
    \actable_shift_57[6]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[6]_net_1\, C => 
        \actable_shift[7]_net_1\, D => refresh, Y => 
        \actable_shift_57[6]_net_1\);
    
    \actable_shift_57_m2[1]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[2]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[1]_net_1\);
    
    \pcable_shift[8]\ : SLE
      port map(D => \pcable_shift_0_sqmuxa_i\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pcable_shift[8]_net_1\);
    
    \rw_p.rwable_shift_7[0]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[1]_net_1\, Y => \rwable_shift_7[0]\);
    
    \rc_shift[5]\ : SLE
      port map(D => \rc_shift_30[5]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[5]_net_1\);
    
    \rc_shift_30[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[6]_net_1\, Y => 
        \rc_shift_30[5]_net_1\);
    
    \pcable_shift[6]\ : SLE
      port map(D => N_765_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \pcable_shift[6]_net_1\);
    
    un1_goactive_4_1 : CFG4
      generic map(INIT => x"0031")

      port map(A => act, B => goact_0, C => \active_0\, D => mode, 
        Y => \un1_goactive_4_1\);
    
    \line[8]\ : SLE
      port map(D => raddr(18), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(8));
    
    active_int : SLE
      port map(D => goact_0, CLK => clk, EN => un36_dopch, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \active_0\);
    
    \actable_shift_57_m2[9]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[10]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[9]_net_1\);
    
    \rw_p.rwable_shift_7[3]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => goact_0, B => un5_dopch_i, C => 
        \rwable_shift[4]_net_1\, Y => \rwable_shift_7[3]\);
    
    \line[0]\ : SLE
      port map(D => raddr(10), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(0));
    
    \rwable_shift[1]\ : SLE
      port map(D => \rwable_shift_7[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[1]_net_1\);
    
    un1_pcable_shift_3_sqmuxa_i_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => bcount(2), B => dorw_0, Y => N_772);
    
    actable_6_iv : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \actable_1_sqmuxa_2\, B => un1_goactive_4_i, 
        C => \actable_shift[0]_net_1\, D => \rc_shift[0]_net_1\, 
        Y => actable_6);
    
    \rc_shift[2]\ : SLE
      port map(D => \rc_shift_30[2]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rc_shift[2]_net_1\);
    
    \line[7]\ : SLE
      port map(D => raddr(17), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(7));
    
    \actable_shift_57[9]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[9]_net_1\, C => 
        \actable_shift[10]_net_1\, D => refresh, Y => 
        \actable_shift_57[9]_net_1\);
    
    \actable_shift_57[11]\ : CFG4
      generic map(INIT => x"F0EE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[11]_net_1\, C => 
        \actable_shift[12]_net_1\, D => refresh, Y => 
        \actable_shift_57[11]_net_1\);
    
    \rc_shift_30[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => goact_0, B => \rc_shift[7]_net_1\, Y => 
        \rc_shift_30[6]_net_1\);
    
    \actable_shift_57[2]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[2]_net_1\, Y => 
        \actable_shift_57[2]_net_1\);
    
    \actable_shift_57[12]\ : CFG4
      generic map(INIT => x"0FEE")

      port map(A => un5_dopch_i, B => 
        \actable_shift_57_m2[12]_net_1\, C => \active_0\, D => 
        refresh, Y => \actable_shift_57[12]_net_1\);
    
    \actable_shift[6]\ : SLE
      port map(D => \actable_shift_57[6]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[6]_net_1\);
    
    un7_dopch : CFG2
      generic map(INIT => x"E")

      port map(A => un5_dopch_i, B => goact_0, Y => un36_dopch);
    
    \pcable_shift_RNO[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => \pcable_shift[4]_net_1\, B => dorw_0, C => 
        bcount(2), Y => N_767_i);
    
    un1_goactive_4 : CFG3
      generic map(INIT => x"10")

      port map(A => refresh, B => un5_dopch_i, C => 
        \un1_goactive_4_1\, Y => un1_goactive_4_i);
    
    actable_shift_57_m2s2 : CFG4
      generic map(INIT => x"FF02")

      port map(A => act, B => goact_0, C => \active_0\, D => mode, 
        Y => actable_shift_57_sm0);
    
    \rwable_shift[0]\ : SLE
      port map(D => \rwable_shift_7[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[0]_net_1\);
    
    \actable_shift_57_m2[2]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[3]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[2]_net_1\);
    
    \rwable_shift[3]\ : SLE
      port map(D => \rwable_shift_7[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rwable_shift[3]_net_1\);
    
    pcable_shift_0_sqmuxa_i : CFG4
      generic map(INIT => x"7FFF")

      port map(A => bcount(1), B => bcount(2), C => dorw_0, D => 
        bcount(0), Y => \pcable_shift_0_sqmuxa_i\);
    
    \actable_shift_57_m2[5]\ : CFG3
      generic map(INIT => x"A8")

      port map(A => \actable_shift[6]_net_1\, B => 
        actable_shift_57_sm0, C => un1_goactive_4_i, Y => 
        \actable_shift_57_m2[5]_net_1\);
    
    \actable_shift[2]\ : SLE
      port map(D => \actable_shift_57[2]_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \actable_shift[2]_net_1\);
    
    \actable_shift_57[5]\ : CFG3
      generic map(INIT => x"54")

      port map(A => refresh, B => un5_dopch_i, C => 
        \actable_shift_57_m2[5]_net_1\, Y => 
        \actable_shift_57[5]_net_1\);
    
    \line[6]\ : SLE
      port map(D => raddr(16), CLK => clk, EN => goact_0, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => line_i_0(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity fastsdram is

    port( raddr           : in    std_logic_vector(30 downto 0);
          b_size          : in    std_logic_vector(3 downto 0);
          ras             : in    std_logic_vector(3 downto 0);
          rcd             : in    std_logic_vector(2 downto 0);
          rrd             : in    std_logic_vector(1 downto 0);
          rp              : in    std_logic_vector(2 downto 0);
          rc              : in    std_logic_vector(3 downto 0);
          rfc             : in    std_logic_vector(3 downto 0);
          wr              : in    std_logic_vector(1 downto 0);
          mrd             : in    std_logic_vector(2 downto 0);
          cl              : in    std_logic_vector(2 downto 0);
          bl              : in    std_logic_vector(1 downto 0);
          ds              : in    std_logic_vector(1 downto 0);
          colbits         : in    std_logic_vector(2 downto 0);
          rowbits         : in    std_logic_vector(1 downto 0);
          sa              : out   std_logic_vector(13 downto 0);
          ba              : out   std_logic_vector(1 downto 0);
          cs_n            : out   std_logic_vector(0 to 0);
          clk             : in    std_logic;
          reset_n         : in    std_logic;
          sd_init         : in    std_logic;
          r_req           : in    std_logic;
          w_req           : in    std_logic;
          auto_pch        : in    std_logic;
          rf_req          : in    std_logic;
          p_req           : in    std_logic;
          m_req           : in    std_logic;
          m_req_dll_reset : in    std_logic;
          em_req          : in    std_logic;
          cl_half         : in    std_logic;
          regdimm         : in    std_logic;
          dqm_wr_bterm    : out   std_logic;
          rw_ack          : out   std_logic;
          s_ack           : out   std_logic;
          r_valid         : out   std_logic;
          w_valid         : out   std_logic;
          d_req           : out   std_logic;
          oe              : out   std_logic;
          cke             : out   std_logic;
          ras_n           : out   std_logic;
          cas_n           : out   std_logic;
          we_n            : out   std_logic
        );

end fastsdram;

architecture DEF_ARCH of fastsdram is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component openbank
    port( wshift_13               : out   std_logic_vector(6 downto 1);
          wshift                  : in    std_logic_vector(6 downto 1) := (others => 'U');
          raddr                   : in    std_logic_vector(22 downto 0) := (others => 'U');
          lnht_cmd                : in    std_logic_vector(3 downto 0) := (others => 'U');
          pcable                  : inout   std_logic_vector(3 downto 0);
          active                  : inout   std_logic_vector(3 downto 0);
          bdcnt                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          rdwr_cmd                : in    std_logic_vector(3 downto 0) := (others => 'U');
          dorw                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          rshift                  : in    std_logic_vector(6 downto 5) := (others => 'U');
          bcount                  : in    std_logic_vector(2 downto 0) := (others => 'U');
          line_i_2                : out   std_logic_vector(11 downto 0);
          bdcnt_6_iv_i_0          : out   std_logic;
          rwable_1                : in    std_logic := 'U';
          rwable_0                : in    std_logic := 'U';
          rwable_3                : in    std_logic := 'U';
          bdcnt_6_2               : out   std_logic;
          bdcnt_6_0               : out   std_logic;
          bdcnt_6_3               : out   std_logic;
          actable_2               : out   std_logic;
          actable_3               : in    std_logic := 'U';
          actable_0               : in    std_logic := 'U';
          cs_n_5_0                : out   std_logic;
          sa_5_5                  : out   std_logic;
          sa_5_1                  : out   std_logic;
          sa_5_0                  : out   std_logic;
          sa_5_10                 : out   std_logic;
          sa_5_8                  : out   std_logic;
          sa_5_2                  : out   std_logic;
          sa_5_3                  : out   std_logic;
          sa_5_4                  : out   std_logic;
          psa_0                   : in    std_logic := 'U';
          psa_8                   : in    std_logic := 'U';
          prch_0                  : in    std_logic := 'U';
          goact_2                 : in    std_logic := 'U';
          goact_0                 : in    std_logic := 'U';
          goact_3                 : in    std_logic := 'U';
          rshift_46_0             : out   std_logic;
          chip_i_2_0              : out   std_logic;
          rw_4                    : out   std_logic;
          N_117_i                 : out   std_logic;
          N_78_i                  : out   std_logic;
          un155_rdwr_cmd          : out   std_logic;
          un197_rdwr_cmd          : out   std_logic;
          un71_rdwr_cmd           : out   std_logic;
          un113_rdwr_cmd          : out   std_logic;
          pchaddr_3_sqmuxa_i_0    : out   std_logic;
          act_4                   : out   std_logic;
          un30_rdwr_cmd           : in    std_logic := 'U';
          un42_rdwr_cmd           : in    std_logic := 'U';
          N_783_i                 : out   std_logic;
          N_77                    : out   std_logic;
          oe_2                    : out   std_logic;
          w_valid_i               : in    std_logic := 'U';
          rc_zero_0_sqmuxa        : out   std_logic;
          wc_zero_0_sqmuxa        : out   std_logic;
          N_812                   : in    std_logic := 'U';
          un222_rdwr_cmd          : out   std_logic;
          un180_rdwr_cmd          : out   std_logic;
          un18_rdwr_cmd           : out   std_logic;
          un54_rdwr_cmd           : out   std_logic;
          un138_rdwr_cmd          : out   std_logic;
          un7_mode_cmd            : out   std_logic;
          un13_rfsh_cmd           : out   std_logic;
          N_73                    : in    std_logic := 'U';
          un13_rfsh_cmd_1         : in    std_logic := 'U';
          we_n_2                  : out   std_logic;
          un16_act_i              : in    std_logic := 'U';
          un1_pch_3_i             : out   std_logic;
          un96_rdwr_cmd           : out   std_logic;
          un1_cs_n_0_sqmuxa_i_0   : in    std_logic := 'U';
          bdzero_2                : out   std_logic;
          bterm_3                 : out   std_logic;
          w_valid_i_1             : out   std_logic;
          rcount_2_sqmuxa         : out   std_logic;
          un217_rdwr_cmd          : out   std_logic;
          turnaround_hold         : in    std_logic := 'U';
          rc_zero_d               : in    std_logic := 'U';
          un1_mode_cmd            : out   std_logic;
          mode_cmd                : in    std_logic := 'U';
          refresh                 : in    std_logic := 'U';
          un4_p_req_0_49_a2_0_a2  : out   std_logic;
          p_req                   : in    std_logic := 'U';
          un1_pch_4_1             : out   std_logic;
          bterm                   : in    std_logic := 'U';
          pchaddr_9_sn_m2_i_1     : out   std_logic;
          pchaddr_9_sn_m3_i_1     : out   std_logic;
          mode                    : in    std_logic := 'U';
          read_cmd                : in    std_logic := 'U';
          un4_rf_req_0_60_a2_0_a2 : out   std_logic;
          rf_req                  : in    std_logic := 'U';
          precharge               : in    std_logic := 'U';
          doread                  : in    std_logic := 'U';
          un36_rw_i_0             : out   std_logic;
          un13_prch_cmd           : out   std_logic;
          rfsh_cmd                : in    std_logic := 'U';
          prch_cmd                : in    std_logic := 'U';
          bdzero                  : in    std_logic := 'U';
          un14_rw                 : in    std_logic := 'U';
          N_125                   : out   std_logic;
          bterm_cmd               : in    std_logic := 'U';
          ack                     : in    std_logic := 'U';
          lnht_cmd26              : out   std_logic;
          un1_rowaddr_int_0_N_2   : in    std_logic := 'U';
          lnht_cmd5               : out   std_logic;
          un1_line_i_0_0_N_2      : in    std_logic := 'U';
          cke                     : in    std_logic := 'U';
          un8_rc_zero             : out   std_logic;
          rc_zero                 : in    std_logic := 'U';
          un4_wc_zero             : out   std_logic;
          wc_zero                 : in    std_logic := 'U';
          dowrite                 : in    std_logic := 'U';
          rw                      : in    std_logic := 'U';
          sa_5_sn_N_4_mux         : in    std_logic := 'U';
          N_6                     : in    std_logic := 'U';
          un78_rw                 : in    std_logic := 'U';
          un1_rw_11_i             : out   std_logic;
          pch                     : in    std_logic := 'U';
          un8_precharge           : in    std_logic := 'U';
          act                     : in    std_logic := 'U';
          clk                     : in    std_logic := 'U';
          reset_n                 : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component openbank_2
    port( bcount     : in    std_logic_vector(2 downto 0) := (others => 'U');
          raddr      : in    std_logic_vector(22 downto 10) := (others => 'U');
          line_i_3   : out   std_logic_vector(11 downto 0);
          prch_0     : in    std_logic := 'U';
          dorw_0     : in    std_logic := 'U';
          actable_0  : out   std_logic;
          rwable_0   : out   std_logic;
          pcable_0   : out   std_logic;
          chip_i_3_0 : out   std_logic;
          active_0   : out   std_logic;
          goact_0    : in    std_logic := 'U';
          refresh    : in    std_logic := 'U';
          mode       : in    std_logic := 'U';
          act        : in    std_logic := 'U';
          read_cmd   : in    std_logic := 'U';
          precharge  : in    std_logic := 'U';
          cke        : in    std_logic := 'U';
          clk        : in    std_logic := 'U';
          reset_n    : in    std_logic := 'U'
        );
  end component;

  component openbank_0
    port( bcount              : in    std_logic_vector(2 downto 0) := (others => 'U');
          raddr               : in    std_logic_vector(22 downto 10) := (others => 'U');
          line_i_1            : out   std_logic_vector(11 downto 0);
          sa_5_0              : out   std_logic;
          sa_5_2              : out   std_logic;
          prch_0              : in    std_logic := 'U';
          dorw_0              : in    std_logic := 'U';
          actable_0           : out   std_logic;
          rwable_0            : out   std_logic;
          pcable_0            : out   std_logic;
          chip_i_1_0          : out   std_logic;
          active_0            : out   std_logic;
          goact_0             : in    std_logic := 'U';
          pch                 : in    std_logic := 'U';
          un8_precharge       : in    std_logic := 'U';
          act                 : in    std_logic := 'U';
          read_cmd            : in    std_logic := 'U';
          precharge           : in    std_logic := 'U';
          cas_n_1             : out   std_logic;
          un1_precharge_5_i_0 : in    std_logic := 'U';
          ras_n_1             : out   std_logic;
          un1_precharge_3_i_0 : in    std_logic := 'U';
          cke                 : in    std_logic := 'U';
          mode                : in    std_logic := 'U';
          refresh             : in    std_logic := 'U';
          clk                 : in    std_logic := 'U';
          reset_n             : in    std_logic := 'U'
        );
  end component;

  component openbank_1
    port( bcount     : in    std_logic_vector(2 downto 0) := (others => 'U');
          raddr      : in    std_logic_vector(22 downto 10) := (others => 'U');
          line_i_0   : out   std_logic_vector(11 downto 0);
          prch_0     : in    std_logic := 'U';
          dorw_0     : in    std_logic := 'U';
          actable_0  : out   std_logic;
          rwable_0   : out   std_logic;
          pcable_0   : out   std_logic;
          chip_i_0_0 : out   std_logic;
          active_0   : out   std_logic;
          goact_0    : in    std_logic := 'U';
          refresh    : in    std_logic := 'U';
          mode       : in    std_logic := 'U';
          act        : in    std_logic := 'U';
          read_cmd   : in    std_logic := 'U';
          precharge  : in    std_logic := 'U';
          cke        : in    std_logic := 'U';
          clk        : in    std_logic := 'U';
          reset_n    : in    std_logic := 'U'
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal cke_net_1, un1_mode_cmd, \goact[2]_net_1\, 
        \dorw[2]_net_1\, \read_cmd\, \prch[2]_net_1\, 
        \actable[2]\, \pcable[2]\, \active[2]\, \line_i_2[0]\, 
        \line_i_2[1]\, \line_i_2[2]\, \line_i_2[3]\, 
        \line_i_2[4]\, \line_i_2[5]\, \line_i_2[6]\, 
        \line_i_2[7]\, \line_i_2[8]\, \line_i_2[9]\, 
        \line_i_2[10]\, \line_i_2[11]\, \chip_i_2[0]\, 
        \goact[1]_net_1\, \dorw[1]_net_1\, \prch[1]_net_1\, 
        \actable[1]\, \rwable[1]\, \pcable[1]\, \active[1]\, 
        \line_i_1[0]\, \line_i_1[1]\, \line_i_1[2]\, 
        \line_i_1[3]\, \line_i_1[4]\, \line_i_1[5]\, 
        \line_i_1[6]\, \line_i_1[7]\, \line_i_1[8]\, 
        \line_i_1[9]\, \line_i_1[10]\, \line_i_1[11]\, 
        \chip_i_1[0]\, \goact[0]_net_1\, \dorw[0]_net_1\, 
        \prch[0]_net_1\, \actable[0]\, \rwable[0]\, \pcable[0]\, 
        \active[0]\, \line_i_0[0]\, \line_i_0[1]\, \line_i_0[2]\, 
        \line_i_0[3]\, \line_i_0[4]\, \line_i_0[5]\, 
        \line_i_0[6]\, \line_i_0[7]\, \line_i_0[8]\, 
        \line_i_0[9]\, \line_i_0[10]\, \line_i_0[11]\, 
        \chip_i_0[0]\, \goact[3]_net_1\, \dorw[3]_net_1\, 
        \prch[3]_net_1\, \actable[3]\, \rwable[3]\, \pcable[3]\, 
        \active[3]\, \line_i_3[0]\, \line_i_3[1]\, \line_i_3[2]\, 
        \line_i_3[3]\, \line_i_3[4]\, \line_i_3[5]\, 
        \line_i_3[6]\, \line_i_3[7]\, \line_i_3[8]\, 
        \line_i_3[9]\, \line_i_3[10]\, \line_i_3[11]\, 
        \chip_i_3[0]\, \wcount[1]_net_1\, \wcount[2]_net_1\, 
        \wcount[3]_net_1\, \rcount[1]_net_1\, \rcount[2]_net_1\, 
        \rcount[3]_net_1\, \bdcnt[2]_net_1\, \bdcnt[3]_net_1\, 
        \oldchip[0]_net_1\, \pchaddr[0]_net_1\, \wc_zero\, 
        \rc_zero\, \lnht_cmd[0]_net_1\, \lnht_cmd[1]_net_1\, 
        \lnht_cmd[2]_net_1\, \lnht_cmd[3]_net_1\, \bterm_cmd\, 
        \ack\, \turnaround_hold\, \bterm\, \prch_cmd\, \rfsh_cmd\, 
        VCC_net_1, \sa[13]\, \dowrite\, \w_valid\, \new_cmd\, 
        \psa_p.un13_prch_cmd\, \dqm_bterm_p.un23_bterm_net_1\, 
        \doread\, \rshift[0]_net_1\, \rc_zero_d\, \mode_cmd\, 
        \psa[8]_net_1\, \bdcnt[0]_net_1\, \bdcnt[1]_net_1\, 
        \act_p.0.un18_rdwr_cmd\, \rdwr_cmd[0]_net_1\, 
        \act_p.1.un30_rdwr_cmd\, \rdwr_cmd[1]_net_1\, 
        \act_p.2.un42_rdwr_cmd\, \rdwr_cmd[2]_net_1\, 
        \act_p.3.un54_rdwr_cmd\, \rdwr_cmd[3]_net_1\, 
        \act_p.0.un96_rdwr_cmd\, \act_p.1.un138_rdwr_cmd\, 
        \act_p.2.un180_rdwr_cmd\, \act_p.3.un217_rdwr_cmd\, 
        \wr_flow_ctrl_p.w_valid_i_1\, \wshift[1]_net_1\, 
        \wcount[0]_net_1\, \act_p.3.un222_rdwr_cmd\, 
        \psa[0]_net_1\, \wr_flow_ctrl_p.oe_2\, 
        \act_p.un13_rfsh_cmd\, \act_p.un7_mode_cmd\, 
        \act_p.act_4\, \act_p.0.un71_rdwr_cmd\, 
        \act_p.1.un113_rdwr_cmd\, \act_p.2.un155_rdwr_cmd\, 
        \act_p.3.un197_rdwr_cmd\, \sd_ctl_p.ba_5[0]_net_1\, 
        \sd_ctl_p.ba_5[1]_net_1\, \cmd_p.un5_r_req\, 
        \act_p.un9_prch_cmd_net_1\, \bterm_p.bterm_3\, 
        \rshift[1]_net_1\, \rshift[2]_net_1\, \rshift[3]_net_1\, 
        \rshift[4]_net_1\, \rshift[5]_net_1\, \rshift[6]_net_1\, 
        \rshift[7]_net_1\, \wshift_13[1]\, \wshift_13[2]\, 
        \wshift_13[3]\, \wshift_13[4]\, \wshift_13[5]\, 
        \wshift_13[6]\, \wshift[2]_net_1\, \wshift[3]_net_1\, 
        \wshift[4]_net_1\, \wshift[5]_net_1\, \wshift[6]_net_1\, 
        \sd_ctl_p.we_n_2\, \act_p.rw_4\, \sd_ctl_p.sa_5[9]\, 
        \sd_ctl_p.sa_5[11]\, \bterm_p.bdzero_2\, 
        \dqs_contention_p.un11_r_req_net_1\, 
        \data_flow_ctrl_p.rshift_46[3]\, 
        \data_flow_ctrl_p.rshift_46[5]\, 
        \data_flow_ctrl_p.rshift_46[6]\, 
        \data_flow_ctrl_p.rshift_46[7]\, \bterm_p.bdcnt_6[0]\, 
        \bterm_p.bdcnt_6[2]\, \bterm_p.bdcnt_6[3]\, 
        \dqs_contention_p.un40_rw_net_1\, \cmd_p.0.lnht_cmd5\, 
        \cmd_p.1.lnht_cmd12_net_1\, \cmd_p.2.lnht_cmd19_net_1\, 
        \cmd_p.3.lnht_cmd26\, \rcount[0]_net_1\, 
        \rc_p.rcount_8[0]\, \rc_p.rcount_8[1]\, 
        \rc_p.rcount_8[2]\, \rc_p.rcount_8[3]\, \mode\, 
        \precharge\, \refresh\, un1_cs_n_0_sqmuxa_i_0, 
        \sd_ctl_p.cs_n_5[0]\, \rw_ack\, \bdzero\, rcount_2_sqmuxa, 
        rc_zero_0_sqmuxa, \rc_p.un8_rc_zero\, un1_precharge_5_i_0, 
        \sd_ctl_p.cas_n_1\, \rc_p.un78_rw_net_1\, 
        wc_zero_0_sqmuxa, \wc_p.un4_wc_zero\, un1_precharge_3_i_0, 
        \sd_ctl_p.ras_n_1\, \bcount[0]_net_1\, \bcount[2]_net_1\, 
        \bcount[1]_net_1\, \bterm_p.op_eq.un14_rw\, un1_rw_11_i, 
        un1_pch_3_i, un16_act_i, un36_rw_i_0, \pch\, 
        \sd_ctl_p.un8_precharge_net_1\, \act\, \sd_ctl_p.sa_5[0]\, 
        \sd_ctl_p.sa_5[1]\, \sd_ctl_p.sa_5[2]\, 
        \sd_ctl_p.sa_5[3]\, \sd_ctl_p.sa_5[4]\, 
        \sd_ctl_p.sa_5[5]\, \sd_ctl_p.sa_5[6]_net_1\, 
        \sd_ctl_p.sa_5[7]_net_1\, \sd_ctl_p.sa_5[8]\, 
        \sd_ctl_p.sa_5[10]\, \mode_cmd_RNO\, 
        \cmd_p.un4_p_req_0_49_a2_0_a2\, 
        \cmd_p.un4_rf_req_0_60_a2_0_a2\, 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_net_1\, 
        \cmd_p.rdwr_cmd_3_1_87_a2_0_a2_net_1\, 
        \cmd_p.rdwr_cmd_3_0_104_a2_0_a2_net_1\, 
        \cmd_p.rdwr_cmd_3_121_a2_0_a2_net_1\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[0]\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[1]\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[2]\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[3]\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[4]\, 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[5]\, 
        \cmd_p.2.un1_rowaddr_int_0_N_2\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[0]\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[1]\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[2]\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[3]\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[4]\, 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[5]\, 
        \cmd_p.1.un1_rowaddr_int_0_N_2\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[0]\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[1]\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[2]\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[3]\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[4]\, 
        \cmd_p.0.un1_line_i_0_0_data_tmp[5]\, 
        \cmd_p.0.un1_line_i_0_0_N_2\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[0]\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[1]\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[2]\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[3]\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[4]\, 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[5]\, 
        \cmd_p.3.un1_rowaddr_int_0_N_2\, pchaddr_3_sqmuxa_i_0, 
        \act_p.un19_rfsh_cmd_net_1\, un1_wc_zero_1_sqmuxa_i, N_74, 
        N_125, \act_p.un13_rfsh_cmd_1\, 
        \act_p.un23_rfsh_cmd_net_1\, \cmd_p.un1_r_req\, 
        \sd_ctl_p.sa_5_sn_N_4_mux\, un1_rcount21, 
        \un16_1.CO1_net_1\, N_73, N_77, N_421, N_422, 
        \rc_p.op_eq.un18_rc_zero\, N_423, N_424, N_812, N_808, 
        \rshift_cnst_7_2_.N_6\, N_56, N_802, N_813, N_798, N_40_i, 
        \act_p.pchaddr_9[0]\, 
        \rc_p.un83_rw_1.un1_wc_zero_1_sqmuxa_i_a3_0_1_net_1\, 
        \openbank_gen.2.openbank_r1_i.un1_pch_4_1\, 
        un1_cs_n_0_sqmuxa_0, \act_p.un23_rfsh_cmd_4_net_1\, 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m2_i_1\, 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m3_i_1\, 
        \rc_p.un72_rw_1.un1_rcount21_0_0_net_1\, \un1_bterm_4_1\, 
        \un1_precharge_5_1\, 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_a3_1_0[7]_net_1\, 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_2[3]_net_1\, 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_0[3]_net_1\, 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_i_0[4]_net_1\, 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\, read_cmd_i, 
        N_117_i, N_78_i, N_783_i, un1_rc_zero_1_sqmuxa_i, N_116_i, 
        N_795_i, N_796_i, N_797_i, \bterm_p.bdcnt_6_iv_i[1]\, 
        N_791_i, N_792_i, N_793_i, N_794_i, 
        \act_p.pchaddr_9_am[0]_net_1\, 
        \act_p.pchaddr_9_ns_1[0]_net_1\, 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns_1[2]_net_1\, 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_1[6]_net_1\, 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_2_1_0[3]_net_1\, 
        \rc_p.un83_rw_1.N_796_i_1_net_1\ : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : openbank
	Use entity work.openbank(DEF_ARCH);
    for all : openbank_2
	Use entity work.openbank_2(DEF_ARCH);
    for all : openbank_0
	Use entity work.openbank_0(DEF_ARCH);
    for all : openbank_1
	Use entity work.openbank_1(DEF_ARCH);
begin 

    sa(13) <= \sa[13]\;
    sa(12) <= \sa[13]\;
    rw_ack <= \rw_ack\;
    w_valid <= \w_valid\;
    d_req <= \sa[13]\;
    cke <= cke_net_1;

    mode_cmd_RNO : CFG4
      generic map(INIT => x"0004")

      port map(A => rf_req, B => m_req, C => \ack\, D => p_req, Y
         => \mode_cmd_RNO\);
    
    \act_p.un23_rfsh_cmd_4\ : CFG2
      generic map(INIT => x"4")

      port map(A => \bterm_cmd\, B => \rfsh_cmd\, Y => 
        \act_p.un13_rfsh_cmd_1\);
    
    \wshift[3]\ : SLE
      port map(D => \wshift_13[3]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[3]_net_1\);
    
    \rshift[3]\ : SLE
      port map(D => \data_flow_ctrl_p.rshift_46[3]\, CLK => clk, 
        EN => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rshift[3]_net_1\);
    
    \ba[0]\ : SLE
      port map(D => \sd_ctl_p.ba_5[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => ba(0));
    
    \rshift[0]\ : SLE
      port map(D => \rshift[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rshift[0]_net_1\);
    
    rc_zero : SLE
      port map(D => un1_rc_zero_1_sqmuxa_i, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rc_zero\);
    
    \cmd_p.2.un1_rowaddr_int_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(13), B => \line_i_2[2]\, C => 
        \line_i_2[3]\, D => raddr(12), FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[1]\);
    
    \dqs_contention_p.un11_r_req\ : CFG4
      generic map(INIT => x"4800")

      port map(A => \oldchip[0]_net_1\, B => \new_cmd\, C => 
        raddr(22), D => r_req, Y => 
        \dqs_contention_p.un11_r_req_net_1\);
    
    \rcount[1]\ : SLE
      port map(D => \rc_p.rcount_8[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rcount[1]_net_1\);
    
    \act_p.1.un30_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \rdwr_cmd[1]_net_1\, B => \actable[1]\, C => 
        N_125, D => \goact[1]_net_1\, Y => 
        \act_p.1.un30_rdwr_cmd\);
    
    ack : SLE
      port map(D => N_117_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \ack\);
    
    pch : SLE
      port map(D => pchaddr_3_sqmuxa_i_0, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => \pch\);
    
    bterm : SLE
      port map(D => \bterm_p.bterm_3\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => \bterm\);
    
    \lnht_cmd[2]\ : SLE
      port map(D => \cmd_p.2.lnht_cmd19_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \lnht_cmd[2]_net_1\);
    
    \sa[5]\ : SLE
      port map(D => \sd_ctl_p.sa_5[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(5));
    
    rw : SLE
      port map(D => \act_p.rw_4\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \rw_ack\);
    
    doread : SLE
      port map(D => \read_cmd\, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \doread\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns_1[2]\ : CFG4
      generic map(INIT => x"4774")

      port map(A => N_798, B => \wc_p.un4_wc_zero\, C => 
        \bcount[1]_net_1\, D => \bcount[2]_net_1\, Y => 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns_1[2]_net_1\);
    
    \bcount[1]\ : SLE
      port map(D => b_size(1), CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \bcount[1]_net_1\);
    
    \wcount[2]\ : SLE
      port map(D => N_792_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \wcount[2]_net_1\);
    
    \un16_1.CO1\ : CFG3
      generic map(INIT => x"F2")

      port map(A => N_421, B => rc_zero_0_sqmuxa, C => N_422, Y
         => \un16_1.CO1_net_1\);
    
    \cmd_p.0.un1_line_i_0_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(13), B => \line_i_0[2]\, C => 
        \line_i_0[3]\, D => raddr(12), FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[1]\);
    
    mode_cmd : SLE
      port map(D => \mode_cmd_RNO\, CLK => clk, EN => N_116_i, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \mode_cmd\);
    
    \bdcnt[3]\ : SLE
      port map(D => \bterm_p.bdcnt_6[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \bdcnt[3]_net_1\);
    
    \rdwr_cmd[3]\ : SLE
      port map(D => \cmd_p.rdwr_cmd_3_121_a2_0_a2_net_1\, CLK => 
        clk, EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rdwr_cmd[3]_net_1\);
    
    \dqm_wr_bterm\ : SLE
      port map(D => \dqm_bterm_p.un23_bterm_net_1\, CLK => clk, 
        EN => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        dqm_wr_bterm);
    
    \we_n\ : SLE
      port map(D => \sd_ctl_p.we_n_2\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => we_n);
    
    \rshift_cnst_7_2_.m1_0_a2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \bcount[2]_net_1\, B => \bcount[1]_net_1\, Y
         => \bterm_p.op_eq.un14_rw\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(15), B => \line_i_3[4]\, C => 
        \line_i_3[5]\, D => raddr(14), FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[2]\);
    
    \rc_p.un72_rw_1.un1_mode_cmd_1[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rc_p.un8_rc_zero\, B => \rcount[2]_net_1\, C
         => \bcount[2]_net_1\, Y => N_423);
    
    \bdcnt[0]\ : SLE
      port map(D => \bterm_p.bdcnt_6[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \bdcnt[0]_net_1\);
    
    \bdcnt[1]\ : SLE
      port map(D => \bterm_p.bdcnt_6_iv_i[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \bdcnt[1]_net_1\);
    
    \ba[1]\ : SLE
      port map(D => \sd_ctl_p.ba_5[1]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => ba(1));
    
    \rdwr_cmd[1]\ : SLE
      port map(D => \cmd_p.rdwr_cmd_3_1_87_a2_0_a2_net_1\, CLK
         => clk, EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rdwr_cmd[1]_net_1\);
    
    \goact[2]\ : SLE
      port map(D => \act_p.2.un42_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \goact[2]_net_1\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0[3]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \rshift[3]_net_1\, B => \rc_p.un78_rw_net_1\, 
        C => un1_rw_11_i, D => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_0[3]_net_1\, 
        Y => \data_flow_ctrl_p.rshift_46[3]\);
    
    \cmd_p.2.un1_rowaddr_int_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(21), B => \line_i_2[10]\, C => 
        \line_i_2[11]\, D => raddr(20), FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[5]\);
    
    \cmd_p.rdwr_cmd_3_1_87_a2_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => raddr(8), B => raddr(9), C => 
        \cmd_p.un1_r_req\, D => 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\, Y => 
        \cmd_p.rdwr_cmd_3_1_87_a2_0_a2_net_1\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(13), B => \line_i_1[2]\, C => 
        \line_i_1[3]\, D => raddr(12), FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[1]\);
    
    \oe\ : SLE
      port map(D => \wr_flow_ctrl_p.oe_2\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => oe);
    
    \dorw[1]\ : SLE
      port map(D => \act_p.1.un113_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \dorw[1]_net_1\);
    
    un1_precharge_5 : CFG4
      generic map(INIT => x"EEFE")

      port map(A => un1_pch_3_i, B => \un1_precharge_5_1\, C => 
        \un1_bterm_4_1\, D => un36_rw_i_0, Y => 
        un1_precharge_5_i_0);
    
    \GND\ : GND
      port map(Y => \sa[13]\);
    
    \rdwr_cmd[0]\ : SLE
      port map(D => \cmd_p.rdwr_cmd_3_0_104_a2_0_a2_net_1\, CLK
         => clk, EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rdwr_cmd[0]_net_1\);
    
    \rc_p.un72_rw_1.rc_p.op_eq.un18_rc_zero\ : CFG3
      generic map(INIT => x"01")

      port map(A => \rcount[3]_net_1\, B => \rcount[2]_net_1\, C
         => \rcount[1]_net_1\, Y => \rc_p.op_eq.un18_rc_zero\);
    
    \prch[3]\ : SLE
      port map(D => \act_p.3.un222_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \prch[3]_net_1\);
    
    \cmd_p.0.un1_line_i_0_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(15), B => \line_i_0[4]\, C => 
        \line_i_0[5]\, D => raddr(14), FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[2]\);
    
    \act_p.un9_prch_cmd\ : CFG4
      generic map(INIT => x"FF02")

      port map(A => \prch_cmd\, B => \precharge\, C => N_73, D
         => \act_p.un23_rfsh_cmd_net_1\, Y => 
        \act_p.un9_prch_cmd_net_1\);
    
    w_valid_i : SLE
      port map(D => \wr_flow_ctrl_p.w_valid_i_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \w_valid\);
    
    \openbank_gen.2.openbank_r1_i\ : openbank
      port map(wshift_13(6) => \wshift_13[6]\, wshift_13(5) => 
        \wshift_13[5]\, wshift_13(4) => \wshift_13[4]\, 
        wshift_13(3) => \wshift_13[3]\, wshift_13(2) => 
        \wshift_13[2]\, wshift_13(1) => \wshift_13[1]\, wshift(6)
         => \wshift[6]_net_1\, wshift(5) => \wshift[5]_net_1\, 
        wshift(4) => \wshift[4]_net_1\, wshift(3) => 
        \wshift[3]_net_1\, wshift(2) => \wshift[2]_net_1\, 
        wshift(1) => \wshift[1]_net_1\, raddr(22) => raddr(22), 
        raddr(21) => raddr(21), raddr(20) => raddr(20), raddr(19)
         => raddr(19), raddr(18) => raddr(18), raddr(17) => 
        raddr(17), raddr(16) => raddr(16), raddr(15) => raddr(15), 
        raddr(14) => raddr(14), raddr(13) => raddr(13), raddr(12)
         => raddr(12), raddr(11) => raddr(11), raddr(10) => 
        raddr(10), raddr(9) => nc2, raddr(8) => nc4, raddr(7) => 
        nc3, raddr(6) => nc1, raddr(5) => raddr(5), raddr(4) => 
        raddr(4), raddr(3) => raddr(3), raddr(2) => raddr(2), 
        raddr(1) => raddr(1), raddr(0) => raddr(0), lnht_cmd(3)
         => \lnht_cmd[3]_net_1\, lnht_cmd(2) => 
        \lnht_cmd[2]_net_1\, lnht_cmd(1) => \lnht_cmd[1]_net_1\, 
        lnht_cmd(0) => \lnht_cmd[0]_net_1\, pcable(3) => 
        \pcable[3]\, pcable(2) => \pcable[2]\, pcable(1) => 
        \pcable[1]\, pcable(0) => \pcable[0]\, active(3) => 
        \active[3]\, active(2) => \active[2]\, active(1) => 
        \active[1]\, active(0) => \active[0]\, bdcnt(3) => 
        \bdcnt[3]_net_1\, bdcnt(2) => \bdcnt[2]_net_1\, bdcnt(1)
         => \bdcnt[1]_net_1\, bdcnt(0) => \bdcnt[0]_net_1\, 
        rdwr_cmd(3) => \rdwr_cmd[3]_net_1\, rdwr_cmd(2) => 
        \rdwr_cmd[2]_net_1\, rdwr_cmd(1) => \rdwr_cmd[1]_net_1\, 
        rdwr_cmd(0) => \rdwr_cmd[0]_net_1\, dorw(3) => 
        \dorw[3]_net_1\, dorw(2) => \dorw[2]_net_1\, dorw(1) => 
        \dorw[1]_net_1\, dorw(0) => \dorw[0]_net_1\, rshift(6)
         => \rshift[6]_net_1\, rshift(5) => \rshift[5]_net_1\, 
        bcount(2) => \bcount[2]_net_1\, bcount(1) => 
        \bcount[1]_net_1\, bcount(0) => \bcount[0]_net_1\, 
        line_i_2(11) => \line_i_2[11]\, line_i_2(10) => 
        \line_i_2[10]\, line_i_2(9) => \line_i_2[9]\, line_i_2(8)
         => \line_i_2[8]\, line_i_2(7) => \line_i_2[7]\, 
        line_i_2(6) => \line_i_2[6]\, line_i_2(5) => 
        \line_i_2[5]\, line_i_2(4) => \line_i_2[4]\, line_i_2(3)
         => \line_i_2[3]\, line_i_2(2) => \line_i_2[2]\, 
        line_i_2(1) => \line_i_2[1]\, line_i_2(0) => 
        \line_i_2[0]\, bdcnt_6_iv_i_0 => 
        \bterm_p.bdcnt_6_iv_i[1]\, rwable_1 => \rwable[1]\, 
        rwable_0 => \rwable[0]\, rwable_3 => \rwable[3]\, 
        bdcnt_6_2 => \bterm_p.bdcnt_6[2]\, bdcnt_6_0 => 
        \bterm_p.bdcnt_6[0]\, bdcnt_6_3 => \bterm_p.bdcnt_6[3]\, 
        actable_2 => \actable[2]\, actable_3 => \actable[3]\, 
        actable_0 => \actable[0]\, cs_n_5_0 => 
        \sd_ctl_p.cs_n_5[0]\, sa_5_5 => \sd_ctl_p.sa_5[5]\, 
        sa_5_1 => \sd_ctl_p.sa_5[1]\, sa_5_0 => 
        \sd_ctl_p.sa_5[0]\, sa_5_10 => \sd_ctl_p.sa_5[10]\, 
        sa_5_8 => \sd_ctl_p.sa_5[8]\, sa_5_2 => 
        \sd_ctl_p.sa_5[2]\, sa_5_3 => \sd_ctl_p.sa_5[3]\, sa_5_4
         => \sd_ctl_p.sa_5[4]\, psa_0 => \psa[0]_net_1\, psa_8
         => \psa[8]_net_1\, prch_0 => \prch[2]_net_1\, goact_2
         => \goact[2]_net_1\, goact_0 => \goact[0]_net_1\, 
        goact_3 => \goact[3]_net_1\, rshift_46_0 => 
        \data_flow_ctrl_p.rshift_46[5]\, chip_i_2_0 => 
        \chip_i_2[0]\, rw_4 => \act_p.rw_4\, N_117_i => N_117_i, 
        N_78_i => N_78_i, un155_rdwr_cmd => 
        \act_p.2.un155_rdwr_cmd\, un197_rdwr_cmd => 
        \act_p.3.un197_rdwr_cmd\, un71_rdwr_cmd => 
        \act_p.0.un71_rdwr_cmd\, un113_rdwr_cmd => 
        \act_p.1.un113_rdwr_cmd\, pchaddr_3_sqmuxa_i_0 => 
        pchaddr_3_sqmuxa_i_0, act_4 => \act_p.act_4\, 
        un30_rdwr_cmd => \act_p.1.un30_rdwr_cmd\, un42_rdwr_cmd
         => \act_p.2.un42_rdwr_cmd\, N_783_i => N_783_i, N_77 => 
        N_77, oe_2 => \wr_flow_ctrl_p.oe_2\, w_valid_i => 
        \w_valid\, rc_zero_0_sqmuxa => rc_zero_0_sqmuxa, 
        wc_zero_0_sqmuxa => wc_zero_0_sqmuxa, N_812 => N_812, 
        un222_rdwr_cmd => \act_p.3.un222_rdwr_cmd\, 
        un180_rdwr_cmd => \act_p.2.un180_rdwr_cmd\, un18_rdwr_cmd
         => \act_p.0.un18_rdwr_cmd\, un54_rdwr_cmd => 
        \act_p.3.un54_rdwr_cmd\, un138_rdwr_cmd => 
        \act_p.1.un138_rdwr_cmd\, un7_mode_cmd => 
        \act_p.un7_mode_cmd\, un13_rfsh_cmd => 
        \act_p.un13_rfsh_cmd\, N_73 => N_73, un13_rfsh_cmd_1 => 
        \act_p.un13_rfsh_cmd_1\, we_n_2 => \sd_ctl_p.we_n_2\, 
        un16_act_i => un16_act_i, un1_pch_3_i => un1_pch_3_i, 
        un96_rdwr_cmd => \act_p.0.un96_rdwr_cmd\, 
        un1_cs_n_0_sqmuxa_i_0 => un1_cs_n_0_sqmuxa_i_0, bdzero_2
         => \bterm_p.bdzero_2\, bterm_3 => \bterm_p.bterm_3\, 
        w_valid_i_1 => \wr_flow_ctrl_p.w_valid_i_1\, 
        rcount_2_sqmuxa => rcount_2_sqmuxa, un217_rdwr_cmd => 
        \act_p.3.un217_rdwr_cmd\, turnaround_hold => 
        \turnaround_hold\, rc_zero_d => \rc_zero_d\, un1_mode_cmd
         => un1_mode_cmd, mode_cmd => \mode_cmd\, refresh => 
        \refresh\, un4_p_req_0_49_a2_0_a2 => 
        \cmd_p.un4_p_req_0_49_a2_0_a2\, p_req => p_req, 
        un1_pch_4_1 => \openbank_gen.2.openbank_r1_i.un1_pch_4_1\, 
        bterm => \bterm\, pchaddr_9_sn_m2_i_1 => 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m2_i_1\, 
        pchaddr_9_sn_m3_i_1 => 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m3_i_1\, 
        mode => \mode\, read_cmd => \read_cmd\, 
        un4_rf_req_0_60_a2_0_a2 => 
        \cmd_p.un4_rf_req_0_60_a2_0_a2\, rf_req => rf_req, 
        precharge => \precharge\, doread => \doread\, un36_rw_i_0
         => un36_rw_i_0, un13_prch_cmd => \psa_p.un13_prch_cmd\, 
        rfsh_cmd => \rfsh_cmd\, prch_cmd => \prch_cmd\, bdzero
         => \bdzero\, un14_rw => \bterm_p.op_eq.un14_rw\, N_125
         => N_125, bterm_cmd => \bterm_cmd\, ack => \ack\, 
        lnht_cmd26 => \cmd_p.3.lnht_cmd26\, un1_rowaddr_int_0_N_2
         => \cmd_p.3.un1_rowaddr_int_0_N_2\, lnht_cmd5 => 
        \cmd_p.0.lnht_cmd5\, un1_line_i_0_0_N_2 => 
        \cmd_p.0.un1_line_i_0_0_N_2\, cke => cke_net_1, 
        un8_rc_zero => \rc_p.un8_rc_zero\, rc_zero => \rc_zero\, 
        un4_wc_zero => \wc_p.un4_wc_zero\, wc_zero => \wc_zero\, 
        dowrite => \dowrite\, rw => \rw_ack\, sa_5_sn_N_4_mux => 
        \sd_ctl_p.sa_5_sn_N_4_mux\, N_6 => \rshift_cnst_7_2_.N_6\, 
        un78_rw => \rc_p.un78_rw_net_1\, un1_rw_11_i => 
        un1_rw_11_i, pch => \pch\, un8_precharge => 
        \sd_ctl_p.un8_precharge_net_1\, act => \act\, clk => clk, 
        reset_n => reset_n);
    
    \cmd_p.2.un1_rowaddr_int_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(11), B => \line_i_2[0]\, C => 
        \line_i_2[1]\, D => raddr(10), FCI => \sa[13]\, S => OPEN, 
        Y => OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[0]\);
    
    \lnht_cmd[0]\ : SLE
      port map(D => \cmd_p.0.lnht_cmd5\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \lnht_cmd[0]_net_1\);
    
    \cmd_p.rdwr_cmd_3_0_104_a2_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => raddr(8), B => raddr(9), C => 
        \cmd_p.un1_r_req\, D => 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\, Y => 
        \cmd_p.rdwr_cmd_3_0_104_a2_0_a2_net_1\);
    
    \cmd_p.2.lnht_cmd19\ : CFG2
      generic map(INIT => x"D")

      port map(A => \cmd_p.2.un1_rowaddr_int_0_N_2\, B => 
        \goact[2]_net_1\, Y => \cmd_p.2.lnht_cmd19_net_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_o3[3]\ : CFG4
      generic map(INIT => x"0ACA")

      port map(A => \wc_zero\, B => \dowrite\, C => \rw_ack\, D
         => N_812, Y => N_802);
    
    \cmd_p.0.un1_line_i_0_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(19), B => \line_i_0[8]\, C => 
        \line_i_0[9]\, D => raddr(18), FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[4]\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(17), B => \line_i_3[6]\, C => 
        \line_i_3[7]\, D => raddr(16), FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[3]\);
    
    \sa[7]\ : SLE
      port map(D => \sd_ctl_p.sa_5[7]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(7));
    
    \rc_p.un83_rw_1.un1_wc_zero_1_sqmuxa_i_a3_0_1\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \wcount[3]_net_1\, B => \wcount[1]_net_1\, C
         => \wcount[2]_net_1\, D => \rc_p.un78_rw_net_1\, Y => 
        \rc_p.un83_rw_1.un1_wc_zero_1_sqmuxa_i_a3_0_1_net_1\);
    
    \cmd_p.rdwr_cmd_3_121_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => raddr(8), B => raddr(9), C => 
        \cmd_p.un1_r_req\, D => 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\, Y => 
        \cmd_p.rdwr_cmd_3_121_a2_0_a2_net_1\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(21), B => \line_i_3[10]\, C => 
        \line_i_3[11]\, D => raddr(20), FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[5]\);
    
    \act_p.pchaddr_9_am[0]\ : CFG4
      generic map(INIT => x"FE10")

      port map(A => 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m3_i_1\, 
        B => N_77, C => \chip_i_1[0]\, D => \chip_i_0[0]\, Y => 
        \act_p.pchaddr_9_am[0]_net_1\);
    
    \sd_ctl_p.un8_precharge\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mode\, B => \bterm\, C => \precharge\, Y => 
        \sd_ctl_p.un8_precharge_net_1\);
    
    bterm_cmd : SLE
      port map(D => N_783_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \bterm_cmd\);
    
    \act_p.un23_rfsh_cmd\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \pcable[2]\, B => \pcable[3]\, C => 
        \act_p.un23_rfsh_cmd_4_net_1\, D => 
        \act_p.un13_rfsh_cmd_1\, Y => \act_p.un23_rfsh_cmd_net_1\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(13), B => \line_i_3[2]\, C => 
        \line_i_3[3]\, D => raddr(12), FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[1]\);
    
    un1_cs_n_0_sqmuxa : CFG4
      generic map(INIT => x"FF01")

      port map(A => \bterm\, B => \pch\, C => raddr(22), D => 
        un1_cs_n_0_sqmuxa_0, Y => un1_cs_n_0_sqmuxa_i_0);
    
    \wshift[4]\ : SLE
      port map(D => \wshift_13[4]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[4]_net_1\);
    
    \rshift[4]\ : SLE
      port map(D => N_795_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \rshift[4]_net_1\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_i_0[4]\ : CFG4
      generic map(INIT => x"0533")

      port map(A => \bcount[2]_net_1\, B => \rshift[5]_net_1\, C
         => un1_rw_11_i, D => \rc_p.un78_rw_net_1\, Y => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_i_0[4]_net_1\);
    
    \pchaddr[0]\ : SLE
      port map(D => \act_p.pchaddr_9[0]\, CLK => clk, EN => 
        pchaddr_3_sqmuxa_i_0, ALn => reset_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \pchaddr[0]_net_1\);
    
    new_cmd : SLE
      port map(D => \ack\, CLK => clk, EN => \cmd_p.un5_r_req\, 
        ALn => reset_n, ADn => \sa[13]\, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \new_cmd\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    rfsh_cmd : SLE
      port map(D => \cmd_p.un4_rf_req_0_60_a2_0_a2\, CLK => clk, 
        EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rfsh_cmd\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_a3_1_0[7]\ : 
        CFG3
      generic map(INIT => x"80")

      port map(A => \bcount[0]_net_1\, B => \bcount[1]_net_1\, C
         => \bcount[2]_net_1\, Y => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_a3_1_0[7]_net_1\);
    
    un1_bterm_4_1 : CFG3
      generic map(INIT => x"02")

      port map(A => \bterm\, B => \mode\, C => \rw_ack\, Y => 
        \un1_bterm_4_1\);
    
    dowrite : SLE
      port map(D => read_cmd_i, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \dowrite\);
    
    \wcount[0]\ : SLE
      port map(D => N_794_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \wcount[0]_net_1\);
    
    \rc_p.un72_rw_1.rc_p.op_eq.un18_rc_zero_RNIK8KR\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \rc_p.un8_rc_zero\, B => 
        \rc_p.op_eq.un18_rc_zero\, C => rc_zero_0_sqmuxa, D => 
        rcount_2_sqmuxa, Y => un1_rc_zero_1_sqmuxa_i);
    
    rc_zero_d : SLE
      port map(D => \rc_zero\, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => \sa[13]\, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \rc_zero_d\);
    
    \cmd_p.un5_r_req_0_o2_0\ : CFG3
      generic map(INIT => x"FE")

      port map(A => p_req, B => m_req, C => rf_req, Y => N_74);
    
    \sa[6]\ : SLE
      port map(D => \sd_ctl_p.sa_5[6]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(6));
    
    \sd_ctl_p.ba_5[0]\ : CFG3
      generic map(INIT => x"02")

      port map(A => raddr(8), B => \precharge\, C => \mode\, Y
         => \sd_ctl_p.ba_5[0]_net_1\);
    
    \rshift_cnst_7_2_.m5\ : CFG3
      generic map(INIT => x"1F")

      port map(A => \bcount[0]_net_1\, B => \bcount[1]_net_1\, C
         => \bcount[2]_net_1\, Y => \rshift_cnst_7_2_.N_6\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(19), B => \line_i_3[8]\, C => 
        \line_i_3[9]\, D => raddr(18), FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[4]\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_1[6]\ : CFG4
      generic map(INIT => x"47CF")

      port map(A => \bcount[2]_net_1\, B => \rc_p.un78_rw_net_1\, 
        C => \rshift[7]_net_1\, D => \bcount[1]_net_1\, Y => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_1[6]_net_1\);
    
    \rcount[2]\ : SLE
      port map(D => \rc_p.rcount_8[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rcount[2]_net_1\);
    
    \rc_p.un78_rw\ : CFG2
      generic map(INIT => x"8")

      port map(A => \rw_ack\, B => \doread\, Y => 
        \rc_p.un78_rw_net_1\);
    
    \rc_p.un72_rw_1.rc_p.rcount_8[0]\ : CFG3
      generic map(INIT => x"09")

      port map(A => N_421, B => rc_zero_0_sqmuxa, C => 
        un1_rcount21, Y => \rc_p.rcount_8[0]\);
    
    \rc_p.un72_rw_1.un1_mode_cmd_1[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \rc_p.un8_rc_zero\, B => \rcount[3]_net_1\, Y
         => N_424);
    
    \prch[0]\ : SLE
      port map(D => \act_p.0.un96_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \prch[0]_net_1\);
    
    \bcount[2]\ : SLE
      port map(D => b_size(2), CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \bcount[2]_net_1\);
    
    \sa[9]\ : SLE
      port map(D => \sd_ctl_p.sa_5[9]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(9));
    
    \cke\ : SLE
      port map(D => VCC_net_1, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => cke_net_1);
    
    \sa[11]\ : SLE
      port map(D => \sd_ctl_p.sa_5[11]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(11));
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_x2_RNI6O0L[1]\ : CFG4
      generic map(INIT => x"0035")

      port map(A => \bcount[1]_net_1\, B => N_40_i, C => 
        \wc_p.un4_wc_zero\, D => N_802, Y => N_793_i);
    
    mode : SLE
      port map(D => \act_p.un7_mode_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => \mode\);
    
    \bdcnt[2]\ : SLE
      port map(D => \bterm_p.bdcnt_6[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \bdcnt[2]_net_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_o2_0_RNIL8RO[3]\ : CFG4
      generic map(INIT => x"0D0F")

      port map(A => \wc_p.un4_wc_zero\, B => \wcount[3]_net_1\, C
         => \rc_p.un83_rw_1.wc_p.wcount_5_i_2[3]_net_1\, D => 
        N_808, Y => N_791_i);
    
    \s_ack\ : SLE
      port map(D => N_78_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => s_ack);
    
    \cmd_p.0.un1_line_i_0_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(17), B => \line_i_0[6]\, C => 
        \line_i_0[7]\, D => raddr(16), FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[3]\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_2_1_0[3]\ : CFG4
      generic map(INIT => x"7FFD")

      port map(A => \wc_p.un4_wc_zero\, B => \rc_p.un78_rw_net_1\, 
        C => \wcount[2]_net_1\, D => N_798, Y => 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_2_1_0[3]_net_1\);
    
    \cmd_p.un5_r_req_0\ : CFG4
      generic map(INIT => x"EEEA")

      port map(A => \ack\, B => \new_cmd\, C => \cmd_p.un1_r_req\, 
        D => N_74, Y => \cmd_p.un5_r_req\);
    
    un1_precharge_3 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mode\, B => \precharge\, C => 
        \openbank_gen.2.openbank_r1_i.un1_pch_4_1\, D => \act\, Y
         => un1_precharge_3_i_0);
    
    \sa[2]\ : SLE
      port map(D => \sd_ctl_p.sa_5[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(2));
    
    \rc_p.un72_rw_1.un1_mode_cmd_1[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rc_p.un8_rc_zero\, B => \rcount[1]_net_1\, C
         => \bcount[1]_net_1\, Y => N_422);
    
    act : SLE
      port map(D => \act_p.act_4\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \act\);
    
    \sa[10]\ : SLE
      port map(D => \sd_ctl_p.sa_5[10]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(10));
    
    \rc_p.un72_rw_1.un1_rcount21_0\ : CFG3
      generic map(INIT => x"DC")

      port map(A => N_812, B => 
        \rc_p.un72_rw_1.un1_rcount21_0_0_net_1\, C => 
        \rc_p.un78_rw_net_1\, Y => un1_rcount21);
    
    \goact[0]\ : SLE
      port map(D => \act_p.0.un18_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \goact[0]_net_1\);
    
    \cmd_p.3.un1_rowaddr_int_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(11), B => \line_i_3[0]\, C => 
        \line_i_3[1]\, D => raddr(10), FCI => \sa[13]\, S => OPEN, 
        Y => OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_data_tmp[0]\);
    
    \wcount[3]\ : SLE
      port map(D => N_791_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \wcount[3]_net_1\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(15), B => \line_i_1[4]\, C => 
        \line_i_1[5]\, D => raddr(14), FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[2]\);
    
    \sd_ctl_p.sa_5[7]\ : CFG4
      generic map(INIT => x"C840")

      port map(A => \act\, B => \sd_ctl_p.sa_5_sn_N_4_mux\, C => 
        raddr(7), D => raddr(17), Y => \sd_ctl_p.sa_5[7]_net_1\);
    
    \psa[8]\ : SLE
      port map(D => \psa_p.un13_prch_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \psa[8]_net_1\);
    
    \dorw[0]\ : SLE
      port map(D => \act_p.0.un71_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \dorw[0]_net_1\);
    
    \openbank_gen.3.openbank_r1_i\ : openbank_2
      port map(bcount(2) => \bcount[2]_net_1\, bcount(1) => 
        \bcount[1]_net_1\, bcount(0) => \bcount[0]_net_1\, 
        raddr(22) => raddr(22), raddr(21) => raddr(21), raddr(20)
         => raddr(20), raddr(19) => raddr(19), raddr(18) => 
        raddr(18), raddr(17) => raddr(17), raddr(16) => raddr(16), 
        raddr(15) => raddr(15), raddr(14) => raddr(14), raddr(13)
         => raddr(13), raddr(12) => raddr(12), raddr(11) => 
        raddr(11), raddr(10) => raddr(10), line_i_3(11) => 
        \line_i_3[11]\, line_i_3(10) => \line_i_3[10]\, 
        line_i_3(9) => \line_i_3[9]\, line_i_3(8) => 
        \line_i_3[8]\, line_i_3(7) => \line_i_3[7]\, line_i_3(6)
         => \line_i_3[6]\, line_i_3(5) => \line_i_3[5]\, 
        line_i_3(4) => \line_i_3[4]\, line_i_3(3) => 
        \line_i_3[3]\, line_i_3(2) => \line_i_3[2]\, line_i_3(1)
         => \line_i_3[1]\, line_i_3(0) => \line_i_3[0]\, prch_0
         => \prch[3]_net_1\, dorw_0 => \dorw[3]_net_1\, actable_0
         => \actable[3]\, rwable_0 => \rwable[3]\, pcable_0 => 
        \pcable[3]\, chip_i_3_0 => \chip_i_3[0]\, active_0 => 
        \active[3]\, goact_0 => \goact[3]_net_1\, refresh => 
        \refresh\, mode => \mode\, act => \act\, read_cmd => 
        \read_cmd\, precharge => \precharge\, cke => cke_net_1, 
        clk => clk, reset_n => reset_n);
    
    \lnht_cmd[3]\ : SLE
      port map(D => \cmd_p.3.lnht_cmd26\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \lnht_cmd[3]_net_1\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_0[3]\ : CFG4
      generic map(INIT => x"0ACC")

      port map(A => N_812, B => \rshift[4]_net_1\, C => 
        un1_rw_11_i, D => \rc_p.un78_rw_net_1\, Y => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_0[3]_net_1\);
    
    \lnht_cmd[1]\ : SLE
      port map(D => \cmd_p.1.lnht_cmd12_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \lnht_cmd[1]_net_1\);
    
    \cmd_p.0.un1_line_i_0_0_I_45\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \chip_i_0[0]\, C => raddr(22), 
        D => \sa[13]\, FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_N_2\);
    
    \rc_p.un72_rw_1.un1_mode_cmd_1[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rc_p.un8_rc_zero\, B => \rcount[0]_net_1\, C
         => \bcount[0]_net_1\, Y => N_421);
    
    \cmd_p.1.lnht_cmd12\ : CFG2
      generic map(INIT => x"D")

      port map(A => \cmd_p.1.un1_rowaddr_int_0_N_2\, B => 
        \goact[1]_net_1\, Y => \cmd_p.1.lnht_cmd12_net_1\);
    
    \sa[0]\ : SLE
      port map(D => \sd_ctl_p.sa_5[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(0));
    
    \cs_n[0]\ : SLE
      port map(D => \sd_ctl_p.cs_n_5[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => cs_n(0));
    
    \act_p.pchaddr_9_ns[0]\ : CFG4
      generic map(INIT => x"4F4A")

      port map(A => \act_p.3.un217_rdwr_cmd\, B => \chip_i_2[0]\, 
        C => \act_p.pchaddr_9_ns_1[0]_net_1\, D => 
        \act_p.pchaddr_9_am[0]_net_1\, Y => \act_p.pchaddr_9[0]\);
    
    \rc_p.un72_rw_1.un1_rcount21_0_0\ : CFG4
      generic map(INIT => x"7340")

      port map(A => \bcount[2]_net_1\, B => \rw_ack\, C => 
        \dowrite\, D => \rc_zero\, Y => 
        \rc_p.un72_rw_1.un1_rcount21_0_0_net_1\);
    
    \cmd_p.0.un1_line_i_0_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(21), B => \line_i_0[10]\, C => 
        \line_i_0[11]\, D => raddr(20), FCI => 
        \cmd_p.0.un1_line_i_0_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[5]\);
    
    \act_p.un5_mode_cmd_i_o2\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \actable[3]\, B => \actable[2]\, C => 
        \actable[1]\, D => \actable[0]\, Y => N_73);
    
    \act_p.un23_rfsh_cmd_4_0\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \precharge\, B => \act_p.un19_rfsh_cmd_net_1\, 
        C => \pcable[0]\, D => \pcable[1]\, Y => 
        \act_p.un23_rfsh_cmd_4_net_1\);
    
    \cmd_p.rdwr_cmd_3_2_71_a2_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => raddr(8), B => raddr(9), C => 
        \cmd_p.un1_r_req\, D => 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\, Y => 
        \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_net_1\);
    
    \rshift[7]\ : SLE
      port map(D => \data_flow_ctrl_p.rshift_46[7]\, CLK => clk, 
        EN => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rshift[7]_net_1\);
    
    \prch[2]\ : SLE
      port map(D => \act_p.2.un180_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \prch[2]_net_1\);
    
    \oldchip[0]\ : SLE
      port map(D => raddr(22), CLK => clk, EN => \rw_ack\, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \oldchip[0]_net_1\);
    
    \rcount[0]\ : SLE
      port map(D => \rc_p.rcount_8[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rcount[0]_net_1\);
    
    \act_p.pchaddr_9_ns_1[0]\ : CFG4
      generic map(INIT => x"3305")

      port map(A => 
        \openbank_gen.2.openbank_r1_i.act_p.pchaddr_9_sn_m2_i_1\, 
        B => \chip_i_3[0]\, C => N_77, D => 
        \act_p.3.un217_rdwr_cmd\, Y => 
        \act_p.pchaddr_9_ns_1[0]_net_1\);
    
    \cas_n\ : SLE
      port map(D => \sd_ctl_p.cas_n_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => cas_n);
    
    \rc_p.un83_rw_1.N_797_i\ : CFG4
      generic map(INIT => x"FA72")

      port map(A => \rc_p.un78_rw_net_1\, B => un1_rw_11_i, C => 
        \rshift[2]_net_1\, D => \rshift[1]_net_1\, Y => N_797_i);
    
    un1_precharge_5_1 : CFG4
      generic map(INIT => x"DDDC")

      port map(A => \mode\, B => \precharge\, C => 
        \openbank_gen.2.openbank_r1_i.un1_pch_4_1\, D => \act\, Y
         => \un1_precharge_5_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_o3_RNI22QN[3]\ : CFG4
      generic map(INIT => x"005C")

      port map(A => \wcount[0]_net_1\, B => \bcount[0]_net_1\, C
         => \wc_p.un4_wc_zero\, D => N_802, Y => N_794_i);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wcount[0]_net_1\, B => \wcount[1]_net_1\, Y
         => N_798);
    
    \bcount[0]\ : SLE
      port map(D => b_size(0), CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \bcount[0]_net_1\);
    
    new_cmd_RNICUUF : CFG2
      generic map(INIT => x"E")

      port map(A => \ack\, B => \new_cmd\, Y => N_116_i);
    
    \prch[1]\ : SLE
      port map(D => \act_p.1.un138_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \prch[1]_net_1\);
    
    \rdwr_cmd[2]\ : SLE
      port map(D => \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_net_1\, CLK
         => clk, EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rdwr_cmd[2]_net_1\);
    
    \rc_p.un83_rw_1.N_796_i_1\ : CFG4
      generic map(INIT => x"47CF")

      port map(A => \bterm_p.op_eq.un14_rw\, B => 
        \rc_p.un78_rw_net_1\, C => \rshift[3]_net_1\, D => 
        \bcount[0]_net_1\, Y => \rc_p.un83_rw_1.N_796_i_1_net_1\);
    
    \rc_p.un72_rw_1.rc_p.rcount_8[3]\ : CFG4
      generic map(INIT => x"00C9")

      port map(A => N_423, B => N_424, C => \un16_1.CO1_net_1\, D
         => un1_rcount21, Y => \rc_p.rcount_8[3]\);
    
    \cmd_p.rdwr_cmd_3_121_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => r_req, B => w_req, Y => \cmd_p.un1_r_req\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_2[3]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \wcount[3]_net_1\, B => N_802, C => 
        \rc_p.un83_rw_1.wc_p.wcount_5_i_2_1_0[3]_net_1\, D => 
        N_56, Y => \rc_p.un83_rw_1.wc_p.wcount_5_i_2[3]_net_1\);
    
    \wshift[6]\ : SLE
      port map(D => \wshift_13[6]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[6]_net_1\);
    
    \rshift[6]\ : SLE
      port map(D => \data_flow_ctrl_p.rshift_46[6]\, CLK => clk, 
        EN => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rshift[6]_net_1\);
    
    \sa[1]\ : SLE
      port map(D => \sd_ctl_p.sa_5[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(1));
    
    \cmd_p.2.un1_rowaddr_int_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(17), B => \line_i_2[6]\, C => 
        \line_i_2[7]\, D => raddr(16), FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[3]\);
    
    \psa[0]\ : SLE
      port map(D => un1_mode_cmd, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \psa[0]_net_1\);
    
    \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => m_req, B => rf_req, C => p_req, D => \ack\, Y
         => \cmd_p.rdwr_cmd_3_2_71_a2_0_a2_0_0_net_1\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(17), B => \line_i_1[6]\, C => 
        \line_i_1[7]\, D => raddr(16), FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[3]\);
    
    \cmd_p.2.un1_rowaddr_int_0_I_45\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \chip_i_2[0]\, C => raddr(22), 
        D => \sa[13]\, FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_N_2\);
    
    \act_p.un19_rfsh_cmd\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \active[2]\, B => \active[1]\, C => 
        \active[3]\, D => \active[0]\, Y => 
        \act_p.un19_rfsh_cmd_net_1\);
    
    \wcount[1]\ : SLE
      port map(D => N_793_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \wcount[1]_net_1\);
    
    un16_act : CFG3
      generic map(INIT => x"10")

      port map(A => \precharge\, B => \mode\, C => \act\, Y => 
        un16_act_i);
    
    \wshift[2]\ : SLE
      port map(D => \wshift_13[2]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[2]_net_1\);
    
    \rshift[2]\ : SLE
      port map(D => N_796_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \rshift[2]_net_1\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0[7]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => \rc_p.un78_rw_net_1\, B => un1_rw_11_i, C => 
        \rshift[7]_net_1\, D => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_a3_1_0[7]_net_1\, 
        Y => \data_flow_ctrl_p.rshift_46[7]\);
    
    \sd_ctl_p.un8_precharge_RNIS0T6\ : CFG2
      generic map(INIT => x"1")

      port map(A => \sd_ctl_p.un8_precharge_net_1\, B => \pch\, Y
         => \sd_ctl_p.sa_5_sn_N_4_mux\);
    
    \goact[3]\ : SLE
      port map(D => \act_p.3.un54_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \goact[3]_net_1\);
    
    \rcount[3]\ : SLE
      port map(D => \rc_p.rcount_8[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rcount[3]_net_1\);
    
    \sa[4]\ : SLE
      port map(D => \sd_ctl_p.sa_5[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(4));
    
    \cmd_p.3.un1_rowaddr_int_0_I_45\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \chip_i_3[0]\, C => raddr(22), 
        D => \sa[13]\, FCI => 
        \cmd_p.3.un1_rowaddr_int_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.3.un1_rowaddr_int_0_N_2\);
    
    \r_valid\ : SLE
      port map(D => \rshift[0]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => r_valid);
    
    turnaround_hold : SLE
      port map(D => \dqs_contention_p.un11_r_req_net_1\, CLK => 
        clk, EN => \dqs_contention_p.un40_rw_net_1\, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \turnaround_hold\);
    
    \openbank_gen.1.openbank_r1_i\ : openbank_0
      port map(bcount(2) => \bcount[2]_net_1\, bcount(1) => 
        \bcount[1]_net_1\, bcount(0) => \bcount[0]_net_1\, 
        raddr(22) => raddr(22), raddr(21) => raddr(21), raddr(20)
         => raddr(20), raddr(19) => raddr(19), raddr(18) => 
        raddr(18), raddr(17) => raddr(17), raddr(16) => raddr(16), 
        raddr(15) => raddr(15), raddr(14) => raddr(14), raddr(13)
         => raddr(13), raddr(12) => raddr(12), raddr(11) => 
        raddr(11), raddr(10) => raddr(10), line_i_1(11) => 
        \line_i_1[11]\, line_i_1(10) => \line_i_1[10]\, 
        line_i_1(9) => \line_i_1[9]\, line_i_1(8) => 
        \line_i_1[8]\, line_i_1(7) => \line_i_1[7]\, line_i_1(6)
         => \line_i_1[6]\, line_i_1(5) => \line_i_1[5]\, 
        line_i_1(4) => \line_i_1[4]\, line_i_1(3) => 
        \line_i_1[3]\, line_i_1(2) => \line_i_1[2]\, line_i_1(1)
         => \line_i_1[1]\, line_i_1(0) => \line_i_1[0]\, sa_5_0
         => \sd_ctl_p.sa_5[9]\, sa_5_2 => \sd_ctl_p.sa_5[11]\, 
        prch_0 => \prch[1]_net_1\, dorw_0 => \dorw[1]_net_1\, 
        actable_0 => \actable[1]\, rwable_0 => \rwable[1]\, 
        pcable_0 => \pcable[1]\, chip_i_1_0 => \chip_i_1[0]\, 
        active_0 => \active[1]\, goact_0 => \goact[1]_net_1\, pch
         => \pch\, un8_precharge => 
        \sd_ctl_p.un8_precharge_net_1\, act => \act\, read_cmd
         => \read_cmd\, precharge => \precharge\, cas_n_1 => 
        \sd_ctl_p.cas_n_1\, un1_precharge_5_i_0 => 
        un1_precharge_5_i_0, ras_n_1 => \sd_ctl_p.ras_n_1\, 
        un1_precharge_3_i_0 => un1_precharge_3_i_0, cke => 
        cke_net_1, mode => \mode\, refresh => \refresh\, clk => 
        clk, reset_n => reset_n);
    
    \cmd_p.2.un1_rowaddr_int_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(15), B => \line_i_2[4]\, C => 
        \line_i_2[5]\, D => raddr(14), FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[2]\);
    
    \rc_p.un72_rw_1.rc_p.rcount_8[1]\ : CFG4
      generic map(INIT => x"0309")

      port map(A => N_421, B => N_422, C => un1_rcount21, D => 
        rc_zero_0_sqmuxa, Y => \rc_p.rcount_8[1]\);
    
    \rc_p.un83_rw_1.un1_wc_zero_1_sqmuxa_i\ : CFG4
      generic map(INIT => x"0F01")

      port map(A => \wc_p.un4_wc_zero\, B => \rc_p.un78_rw_net_1\, 
        C => wc_zero_0_sqmuxa, D => 
        \rc_p.un83_rw_1.un1_wc_zero_1_sqmuxa_i_a3_0_1_net_1\, Y
         => un1_wc_zero_1_sqmuxa_i);
    
    \dqs_contention_p.un40_rw\ : CFG2
      generic map(INIT => x"E")

      port map(A => \dqs_contention_p.un11_r_req_net_1\, B => 
        \rw_ack\, Y => \dqs_contention_p.un40_rw_net_1\);
    
    \sa[3]\ : SLE
      port map(D => \sd_ctl_p.sa_5[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(3));
    
    wc_zero : SLE
      port map(D => un1_wc_zero_1_sqmuxa_i, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \wc_zero\);
    
    precharge : SLE
      port map(D => \act_p.un9_prch_cmd_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \precharge\);
    
    \rc_p.un72_rw_1.rc_p.rcount_8[2]\ : CFG3
      generic map(INIT => x"21")

      port map(A => N_423, B => un1_rcount21, C => 
        \un16_1.CO1_net_1\, Y => \rc_p.rcount_8[2]\);
    
    \cmd_p.2.un1_rowaddr_int_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(19), B => \line_i_2[8]\, C => 
        \line_i_2[9]\, D => raddr(18), FCI => 
        \cmd_p.2.un1_rowaddr_int_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.2.un1_rowaddr_int_0_data_tmp[4]\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(19), B => \line_i_1[8]\, C => 
        \line_i_1[9]\, D => raddr(18), FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[4]\);
    
    \dorw[2]\ : SLE
      port map(D => \act_p.2.un155_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \dorw[2]_net_1\);
    
    \sd_ctl_p.sa_5[6]\ : CFG4
      generic map(INIT => x"C840")

      port map(A => \act\, B => \sd_ctl_p.sa_5_sn_N_4_mux\, C => 
        raddr(6), D => raddr(16), Y => \sd_ctl_p.sa_5[6]_net_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns_RNI7DFH[2]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_813, B => N_802, Y => N_792_i);
    
    \ras_n\ : SLE
      port map(D => \sd_ctl_p.ras_n_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => ras_n);
    
    \dqm_bterm_p.un23_bterm\ : CFG2
      generic map(INIT => x"8")

      port map(A => \bterm\, B => \w_valid\, Y => 
        \dqm_bterm_p.un23_bterm_net_1\);
    
    \openbank_gen.0.openbank_r1_i\ : openbank_1
      port map(bcount(2) => \bcount[2]_net_1\, bcount(1) => 
        \bcount[1]_net_1\, bcount(0) => \bcount[0]_net_1\, 
        raddr(22) => raddr(22), raddr(21) => raddr(21), raddr(20)
         => raddr(20), raddr(19) => raddr(19), raddr(18) => 
        raddr(18), raddr(17) => raddr(17), raddr(16) => raddr(16), 
        raddr(15) => raddr(15), raddr(14) => raddr(14), raddr(13)
         => raddr(13), raddr(12) => raddr(12), raddr(11) => 
        raddr(11), raddr(10) => raddr(10), line_i_0(11) => 
        \line_i_0[11]\, line_i_0(10) => \line_i_0[10]\, 
        line_i_0(9) => \line_i_0[9]\, line_i_0(8) => 
        \line_i_0[8]\, line_i_0(7) => \line_i_0[7]\, line_i_0(6)
         => \line_i_0[6]\, line_i_0(5) => \line_i_0[5]\, 
        line_i_0(4) => \line_i_0[4]\, line_i_0(3) => 
        \line_i_0[3]\, line_i_0(2) => \line_i_0[2]\, line_i_0(1)
         => \line_i_0[1]\, line_i_0(0) => \line_i_0[0]\, prch_0
         => \prch[0]_net_1\, dorw_0 => \dorw[0]_net_1\, actable_0
         => \actable[0]\, rwable_0 => \rwable[0]\, pcable_0 => 
        \pcable[0]\, chip_i_0_0 => \chip_i_0[0]\, active_0 => 
        \active[0]\, goact_0 => \goact[0]_net_1\, refresh => 
        \refresh\, mode => \mode\, act => \act\, read_cmd => 
        \read_cmd\, precharge => \precharge\, cke => cke_net_1, 
        clk => clk, reset_n => reset_n);
    
    bdzero : SLE
      port map(D => \bterm_p.bdzero_2\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => \bdzero\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_a3[3]\ : CFG4
      generic map(INIT => x"007E")

      port map(A => \bcount[2]_net_1\, B => \bcount[1]_net_1\, C
         => \rc_p.un78_rw_net_1\, D => \wc_p.un4_wc_zero\, Y => 
        N_56);
    
    \wshift[1]\ : SLE
      port map(D => \wshift_13[1]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[1]_net_1\);
    
    \rshift[1]\ : SLE
      port map(D => N_797_i, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \rshift[1]_net_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_x2[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wcount[0]_net_1\, B => \wcount[1]_net_1\, Y
         => N_40_i);
    
    \dorw[3]\ : SLE
      port map(D => \act_p.3.un197_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \dorw[3]_net_1\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(11), B => \line_i_1[0]\, C => 
        \line_i_1[1]\, D => raddr(10), FCI => \sa[13]\, S => OPEN, 
        Y => OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[0]\);
    
    \wshift[5]\ : SLE
      port map(D => \wshift_13[5]\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \wshift[5]_net_1\);
    
    \rshift[5]\ : SLE
      port map(D => \data_flow_ctrl_p.rshift_46[5]\, CLK => clk, 
        EN => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \rshift[5]_net_1\);
    
    \sa[8]\ : SLE
      port map(D => \sd_ctl_p.sa_5[8]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => sa(8));
    
    read_cmd : SLE
      port map(D => r_req, CLK => clk, EN => VCC_net_1, ALn => 
        reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \read_cmd\);
    
    \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0[6]\ : CFG4
      generic map(INIT => x"80DF")

      port map(A => \rc_p.un78_rw_net_1\, B => \rshift[6]_net_1\, 
        C => un1_rw_11_i, D => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_0_1[6]_net_1\, 
        Y => \data_flow_ctrl_p.rshift_46[6]\);
    
    \rc_p.un83_rw_1.N_796_i\ : CFG4
      generic map(INIT => x"8AD5")

      port map(A => \rc_p.un78_rw_net_1\, B => \rshift[2]_net_1\, 
        C => un1_rw_11_i, D => \rc_p.un83_rw_1.N_796_i_1_net_1\, 
        Y => N_796_i);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns[2]\ : CFG4
      generic map(INIT => x"2DD2")

      port map(A => \wc_p.un4_wc_zero\, B => \wcount[2]_net_1\, C
         => \rc_p.un83_rw_1.wc_p.wcount_5_i_m3_ns_1[2]_net_1\, D
         => \rc_p.un78_rw_net_1\, Y => N_813);
    
    dowrite_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \read_cmd\, Y => read_cmd_i);
    
    \act_p.2.un42_rdwr_cmd_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \rdwr_cmd[2]_net_1\, B => \actable[2]\, C => 
        N_125, D => \goact[2]_net_1\, Y => 
        \act_p.2.un42_rdwr_cmd\);
    
    refresh : SLE
      port map(D => \act_p.un13_rfsh_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \refresh\);
    
    \goact[1]\ : SLE
      port map(D => \act_p.1.un30_rdwr_cmd\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \goact[1]_net_1\);
    
    \cmd_p.1.un1_rowaddr_int_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(21), B => \line_i_1[10]\, C => 
        \line_i_1[11]\, D => raddr(20), FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_data_tmp[5]\);
    
    \cmd_p.0.un1_line_i_0_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => raddr(11), B => \line_i_0[0]\, C => 
        \line_i_0[1]\, D => raddr(10), FCI => \sa[13]\, S => OPEN, 
        Y => OPEN, FCO => \cmd_p.0.un1_line_i_0_0_data_tmp[0]\);
    
    \rc_p.un83_rw_1.N_795_i\ : CFG4
      generic map(INIT => x"00BF")

      port map(A => \rshift[4]_net_1\, B => \rc_p.un78_rw_net_1\, 
        C => un1_rw_11_i, D => 
        \rc_p.un83_rw_1.data_flow_ctrl_p.rshift_46_i_0[4]_net_1\, 
        Y => N_795_i);
    
    \cmd_p.1.un1_rowaddr_int_0_I_45\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \chip_i_1[0]\, C => raddr(22), 
        D => \sa[13]\, FCI => 
        \cmd_p.1.un1_rowaddr_int_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \cmd_p.1.un1_rowaddr_int_0_N_2\);
    
    un1_cs_n_0_sqmuxa_0_0 : CFG4
      generic map(INIT => x"5530")

      port map(A => \oldchip[0]_net_1\, B => \pchaddr[0]_net_1\, 
        C => \pch\, D => \bterm\, Y => un1_cs_n_0_sqmuxa_0);
    
    \rc_p.un83_rw_1.CO2_i_a2_i_o3\ : CFG3
      generic map(INIT => x"F8")

      port map(A => \bcount[0]_net_1\, B => \bcount[1]_net_1\, C
         => \bcount[2]_net_1\, Y => N_812);
    
    \sd_ctl_p.ba_5[1]\ : CFG3
      generic map(INIT => x"02")

      port map(A => raddr(9), B => \precharge\, C => \mode\, Y
         => \sd_ctl_p.ba_5[1]_net_1\);
    
    \rc_p.un83_rw_1.wc_p.wcount_5_i_o2_0[3]\ : CFG3
      generic map(INIT => x"7E")

      port map(A => \rc_p.un78_rw_net_1\, B => \wcount[2]_net_1\, 
        C => N_798, Y => N_808);
    
    prch_cmd : SLE
      port map(D => \cmd_p.un4_p_req_0_49_a2_0_a2\, CLK => clk, 
        EN => N_116_i, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \prch_cmd\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity fastinit is

    port( raddr    : in    std_logic_vector(30 downto 0);
          b_size   : in    std_logic_vector(3 downto 0);
          ras      : in    std_logic_vector(3 downto 0);
          rcd      : in    std_logic_vector(2 downto 0);
          rrd      : in    std_logic_vector(1 downto 0);
          rp       : in    std_logic_vector(2 downto 0);
          rc       : in    std_logic_vector(3 downto 0);
          rfc      : in    std_logic_vector(3 downto 0);
          wr       : in    std_logic_vector(1 downto 0);
          mrd      : in    std_logic_vector(2 downto 0);
          cl       : in    std_logic_vector(2 downto 0);
          bl       : in    std_logic_vector(1 downto 0);
          ds       : in    std_logic_vector(1 downto 0);
          delay    : in    std_logic_vector(15 downto 0);
          ref      : in    std_logic_vector(15 downto 0);
          colbits  : in    std_logic_vector(2 downto 0);
          rowbits  : in    std_logic_vector(1 downto 0);
          sa       : out   std_logic_vector(13 downto 0);
          ba       : out   std_logic_vector(1 downto 0);
          cs_n     : out   std_logic_vector(0 to 0);
          clk      : in    std_logic;
          reset_n  : in    std_logic;
          r_req    : in    std_logic;
          w_req    : in    std_logic;
          auto_pch : in    std_logic;
          sd_init  : in    std_logic;
          cl_half  : in    std_logic;
          regdimm  : in    std_logic;
          rw_ack   : out   std_logic;
          r_valid  : out   std_logic;
          d_req    : out   std_logic;
          w_valid  : out   std_logic;
          oe       : out   std_logic;
          dqm      : out   std_logic;
          cke      : out   std_logic;
          ras_n    : out   std_logic;
          cas_n    : out   std_logic;
          we_n     : out   std_logic
        );

end fastinit;

architecture DEF_ARCH of fastinit is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component fastsdram
    port( raddr           : in    std_logic_vector(30 downto 0) := (others => 'U');
          b_size          : in    std_logic_vector(3 downto 0) := (others => 'U');
          ras             : in    std_logic_vector(3 downto 0) := (others => 'U');
          rcd             : in    std_logic_vector(2 downto 0) := (others => 'U');
          rrd             : in    std_logic_vector(1 downto 0) := (others => 'U');
          rp              : in    std_logic_vector(2 downto 0) := (others => 'U');
          rc              : in    std_logic_vector(3 downto 0) := (others => 'U');
          rfc             : in    std_logic_vector(3 downto 0) := (others => 'U');
          wr              : in    std_logic_vector(1 downto 0) := (others => 'U');
          mrd             : in    std_logic_vector(2 downto 0) := (others => 'U');
          cl              : in    std_logic_vector(2 downto 0) := (others => 'U');
          bl              : in    std_logic_vector(1 downto 0) := (others => 'U');
          ds              : in    std_logic_vector(1 downto 0) := (others => 'U');
          colbits         : in    std_logic_vector(2 downto 0) := (others => 'U');
          rowbits         : in    std_logic_vector(1 downto 0) := (others => 'U');
          sa              : out   std_logic_vector(13 downto 0);
          ba              : out   std_logic_vector(1 downto 0);
          cs_n            : out   std_logic_vector(0 to 0);
          clk             : in    std_logic := 'U';
          reset_n         : in    std_logic := 'U';
          sd_init         : in    std_logic := 'U';
          r_req           : in    std_logic := 'U';
          w_req           : in    std_logic := 'U';
          auto_pch        : in    std_logic := 'U';
          rf_req          : in    std_logic := 'U';
          p_req           : in    std_logic := 'U';
          m_req           : in    std_logic := 'U';
          m_req_dll_reset : in    std_logic := 'U';
          em_req          : in    std_logic := 'U';
          cl_half         : in    std_logic := 'U';
          regdimm         : in    std_logic := 'U';
          dqm_wr_bterm    : out   std_logic;
          rw_ack          : out   std_logic;
          s_ack           : out   std_logic;
          r_valid         : out   std_logic;
          w_valid         : out   std_logic;
          d_req           : out   std_logic;
          oe              : out   std_logic;
          cke             : out   std_logic;
          ras_n           : out   std_logic;
          cas_n           : out   std_logic;
          we_n            : out   std_logic
        );
  end component;

    signal un4_timer_cry_1_S, un4_timer_cry_2_S, 
        un4_timer_cry_3_S, un4_timer_cry_4_S, un4_timer_cry_5_S, 
        un4_timer_cry_6_S, un4_timer_cry_7_S, un4_timer_cry_8_S, 
        un4_timer_cry_9_S, un4_timer_cry_10_S, un4_timer_cry_11_S, 
        un4_timer_cry_12_S, un4_timer_cry_13_S, 
        un4_timer_cry_14_S, un4_timer_s_15_S, \r_req_i\, 
        \w_req_i\, \rf_req\, \m_req\, \sa[13]\, dqm_wr_bterm, 
        s_ack, \timer[0]_net_1\, \timer[1]_net_1\, 
        \timer[2]_net_1\, \timer[3]_net_1\, \timer[4]_net_1\, 
        \timer[5]_net_1\, \timer[6]_net_1\, \timer[7]_net_1\, 
        \timer[8]_net_1\, \timer[9]_net_1\, \timer[10]_net_1\, 
        \timer[11]_net_1\, \timer[12]_net_1\, \timer[13]_net_1\, 
        \timer[14]_net_1\, \timer[15]_net_1\, \r_shift[9]_net_1\, 
        VCC_net_1, \dqm_init_d0\, \dqm_init\, \start_delay_done\, 
        \dqm_init_p.un6_m_req_net_1\, \dqm_init_d1\, \inited\, 
        \m_shift[0]_net_1\, \r_shift[0]_net_1\, 
        \m_shift[1]_net_1\, \m_shift[2]_net_1\, 
        \m_shift[3]_net_1\, \m_shift[4]_net_1\, 
        \m_shift[5]_net_1\, \m_shift[6]_net_1\, 
        \m_shift[7]_net_1\, p_req, \m_shift[9]_net_1\, 
        \r_shift[1]_net_1\, \r_shift[2]_net_1\, 
        \r_shift[3]_net_1\, \r_shift[4]_net_1\, 
        \r_shift[5]_net_1\, \r_shift[6]_net_1\, 
        \r_shift[7]_net_1\, \r_shift[8]_net_1\, 
        \init.un5_timer_reset_net_1\, 
        \timer_p.timer_reset_2_net_1\, \timer_p.timer_6[0]\, 
        \timer_p.timer_6[1]\, \timer_p.timer_6[2]\, 
        \timer_p.timer_6[3]\, \timer_p.timer_6[4]\, 
        \timer_p.timer_6[5]\, \timer_p.timer_6[6]\, 
        \timer_p.timer_6[7]\, \timer_p.timer_6[8]\, 
        \timer_p.timer_6[9]\, \timer_p.timer_6[10]\, 
        \timer_p.timer_6[11]\, \timer_p.timer_6[12]\, 
        \timer_p.timer_6[13]\, \timer_p.timer_6[14]\, 
        \timer_p.timer_6[15]\, \r_shift_0[9]_net_1\, \load\, 
        \timer_reset\, \un4_timer_cry_0\, \un4_timer_cry_1\, 
        \un4_timer_cry_2\, \un4_timer_cry_3\, \un4_timer_cry_4\, 
        \un4_timer_cry_5\, \un4_timer_cry_6\, \un4_timer_cry_7\, 
        \un4_timer_cry_8\, \un4_timer_cry_9\, \un4_timer_cry_10\, 
        \un4_timer_cry_11\, \un4_timer_cry_12\, 
        \un4_timer_cry_13\, \un4_timer_cry_14\, 
        \timer_p.timer_reset_2_0_net_1\, 
        \timer_p.timer_reset_2_9_net_1\, 
        \timer_p.timer_reset_2_10_net_1\, 
        \timer_p.timer_reset_2_11_net_1\, 
        \timer_p.timer_reset_2_12_net_1\, un1_dll_holdoff_en2_i
         : std_logic;
    signal nc2, nc1 : std_logic;

    for all : fastsdram
	Use entity work.fastsdram(DEF_ARCH);
begin 

    sa(13) <= \sa[13]\;
    sa(12) <= \sa[13]\;
    d_req <= \sa[13]\;

    \timer[6]\ : SLE
      port map(D => \timer_p.timer_6[6]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[6]_net_1\);
    
    \timer_RNO[12]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_12_S, Y => \timer_p.timer_6[12]\);
    
    \timer_p.timer_reset_2_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => \timer[1]_net_1\, B => \timer[15]_net_1\, Y
         => \timer_p.timer_reset_2_0_net_1\);
    
    \timer[11]\ : SLE
      port map(D => \timer_p.timer_6[11]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[11]_net_1\);
    
    \m_shift[0]\ : SLE
      port map(D => \m_shift[1]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[0]_net_1\);
    
    un4_timer_cry_0 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[0]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \sa[13]\, S => OPEN, Y
         => OPEN, FCO => \un4_timer_cry_0\);
    
    \r_shift[2]\ : SLE
      port map(D => \r_shift[3]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[2]_net_1\);
    
    \timer_RNO[5]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_5_S, Y => \timer_p.timer_6[5]\);
    
    \timer[9]\ : SLE
      port map(D => \timer_p.timer_6[9]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[9]_net_1\);
    
    un4_timer_cry_8 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[8]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_7\, S => 
        un4_timer_cry_8_S, Y => OPEN, FCO => \un4_timer_cry_8\);
    
    \r_shift[3]\ : SLE
      port map(D => \r_shift[4]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[3]_net_1\);
    
    \timer_RNO[0]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \load\, B => \timer_reset\, C => 
        \timer[0]_net_1\, Y => \timer_p.timer_6[0]\);
    
    \m_shift[7]\ : SLE
      port map(D => p_req, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[7]_net_1\);
    
    un4_timer_cry_10 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[10]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_9\, S => 
        un4_timer_cry_10_S, Y => OPEN, FCO => \un4_timer_cry_10\);
    
    dqm_init_d1 : SLE
      port map(D => \dqm_init_d0\, CLK => clk, EN => VCC_net_1, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \dqm_init_d1\);
    
    \timer_p.timer_6_f0[11]\ : CFG3
      generic map(INIT => x"32")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_11_S, Y => \timer_p.timer_6[11]\);
    
    un4_timer_cry_14 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[14]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_13\, S => 
        un4_timer_cry_14_S, Y => OPEN, FCO => \un4_timer_cry_14\);
    
    \timer[8]\ : SLE
      port map(D => \timer_p.timer_6[8]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[8]_net_1\);
    
    \timer[2]\ : SLE
      port map(D => \timer_p.timer_6[2]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => \sa[13]\, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[2]_net_1\);
    
    \m_shift[2]\ : SLE
      port map(D => \m_shift[3]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[2]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \timer[4]\ : SLE
      port map(D => \timer_p.timer_6[4]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[4]_net_1\);
    
    un4_timer_cry_13 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[13]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_12\, S => 
        un4_timer_cry_13_S, Y => OPEN, FCO => \un4_timer_cry_13\);
    
    timer_reset : SLE
      port map(D => \timer_p.timer_reset_2_net_1\, CLK => clk, EN
         => VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer_reset\);
    
    \timer_p.timer_reset_2_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \timer[13]_net_1\, B => \timer[12]_net_1\, C
         => \timer[11]_net_1\, D => \timer[10]_net_1\, Y => 
        \timer_p.timer_reset_2_11_net_1\);
    
    \timer[1]\ : SLE
      port map(D => \timer_p.timer_6[1]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[1]_net_1\);
    
    \m_shift[5]\ : SLE
      port map(D => \m_shift[6]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[5]_net_1\);
    
    \r_shift[8]\ : SLE
      port map(D => \r_shift[9]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[8]_net_1\);
    
    \dqm\ : CFG2
      generic map(INIT => x"E")

      port map(A => \dqm_init_d1\, B => dqm_wr_bterm, Y => dqm);
    
    \timer_RNO[1]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_1_S, Y => \timer_p.timer_6[1]\);
    
    m_req : SLE
      port map(D => \m_shift[0]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_req\);
    
    \timer_RNO[13]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_13_S, Y => \timer_p.timer_6[13]\);
    
    \timer[15]\ : SLE
      port map(D => \timer_p.timer_6[15]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[15]_net_1\);
    
    \timer_RNO[6]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_6_S, Y => \timer_p.timer_6[6]\);
    
    \r_shift[9]\ : SLE
      port map(D => \r_shift_0[9]_net_1\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \r_shift[9]_net_1\);
    
    \timer_RNO[10]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_10_S, Y => \timer_p.timer_6[10]\);
    
    \dqm_init_p.un6_m_req\ : CFG2
      generic map(INIT => x"8")

      port map(A => \m_req\, B => s_ack, Y => 
        \dqm_init_p.un6_m_req_net_1\);
    
    load : SLE
      port map(D => \sa[13]\, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => \sa[13]\, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \load\);
    
    \m_shift[3]\ : SLE
      port map(D => \m_shift[4]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[3]_net_1\);
    
    \m_shift[9]\ : SLE
      port map(D => \sa[13]\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[9]_net_1\);
    
    \timer[0]\ : SLE
      port map(D => \timer_p.timer_6[0]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[0]_net_1\);
    
    \GND\ : GND
      port map(Y => \sa[13]\);
    
    un4_timer_cry_4 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[4]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_3\, S => 
        un4_timer_cry_4_S, Y => OPEN, FCO => \un4_timer_cry_4\);
    
    \timer_p.timer_reset_2_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \timer[9]_net_1\, B => \timer[8]_net_1\, C
         => \timer[7]_net_1\, D => \timer[6]_net_1\, Y => 
        \timer_p.timer_reset_2_10_net_1\);
    
    inited : SLE
      port map(D => \dqm_init_p.un6_m_req_net_1\, CLK => clk, EN
         => un1_dll_holdoff_en2_i, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \inited\);
    
    start_delay_done : SLE
      port map(D => VCC_net_1, CLK => clk, EN => \timer_reset\, 
        ALn => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => \sa[13]\, LAT => \sa[13]\, Q => \start_delay_done\);
    
    \timer_RNO[15]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_s_15_S, Y => \timer_p.timer_6[15]\);
    
    \timer[3]\ : SLE
      port map(D => \timer_p.timer_6[3]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[3]_net_1\);
    
    \timer_p.timer_6_f0[9]\ : CFG3
      generic map(INIT => x"32")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_9_S, Y => \timer_p.timer_6[9]\);
    
    un4_timer_cry_5 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[5]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_4\, S => 
        un4_timer_cry_5_S, Y => OPEN, FCO => \un4_timer_cry_5\);
    
    un4_timer_cry_1 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[1]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_0\, S => 
        un4_timer_cry_1_S, Y => OPEN, FCO => \un4_timer_cry_1\);
    
    un4_timer_cry_9 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[9]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_8\, S => 
        un4_timer_cry_9_S, Y => OPEN, FCO => \un4_timer_cry_9\);
    
    un4_timer_cry_6 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[6]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_5\, S => 
        un4_timer_cry_6_S, Y => OPEN, FCO => \un4_timer_cry_6\);
    
    fastsdram_1 : fastsdram
      port map(raddr(30) => \sa[13]\, raddr(29) => \sa[13]\, 
        raddr(28) => \sa[13]\, raddr(27) => \sa[13]\, raddr(26)
         => \sa[13]\, raddr(25) => \sa[13]\, raddr(24) => 
        \sa[13]\, raddr(23) => \sa[13]\, raddr(22) => raddr(22), 
        raddr(21) => raddr(21), raddr(20) => raddr(20), raddr(19)
         => raddr(19), raddr(18) => raddr(18), raddr(17) => 
        raddr(17), raddr(16) => raddr(16), raddr(15) => raddr(15), 
        raddr(14) => raddr(14), raddr(13) => raddr(13), raddr(12)
         => raddr(12), raddr(11) => raddr(11), raddr(10) => 
        raddr(10), raddr(9) => raddr(9), raddr(8) => raddr(8), 
        raddr(7) => raddr(7), raddr(6) => raddr(6), raddr(5) => 
        raddr(5), raddr(4) => raddr(4), raddr(3) => raddr(3), 
        raddr(2) => raddr(2), raddr(1) => raddr(1), raddr(0) => 
        raddr(0), b_size(3) => \sa[13]\, b_size(2) => b_size(2), 
        b_size(1) => b_size(1), b_size(0) => b_size(0), ras(3)
         => \sa[13]\, ras(2) => \sa[13]\, ras(1) => VCC_net_1, 
        ras(0) => \sa[13]\, rcd(2) => \sa[13]\, rcd(1) => 
        VCC_net_1, rcd(0) => \sa[13]\, rrd(1) => VCC_net_1, 
        rrd(0) => \sa[13]\, rp(2) => \sa[13]\, rp(1) => VCC_net_1, 
        rp(0) => VCC_net_1, rc(3) => VCC_net_1, rc(2) => \sa[13]\, 
        rc(1) => \sa[13]\, rc(0) => \sa[13]\, rfc(3) => VCC_net_1, 
        rfc(2) => \sa[13]\, rfc(1) => \sa[13]\, rfc(0) => 
        VCC_net_1, wr(1) => VCC_net_1, wr(0) => \sa[13]\, mrd(2)
         => \sa[13]\, mrd(1) => VCC_net_1, mrd(0) => \sa[13]\, 
        cl(2) => \sa[13]\, cl(1) => VCC_net_1, cl(0) => \sa[13]\, 
        bl(1) => VCC_net_1, bl(0) => VCC_net_1, ds(1) => \sa[13]\, 
        ds(0) => \sa[13]\, colbits(2) => \sa[13]\, colbits(1) => 
        VCC_net_1, colbits(0) => VCC_net_1, rowbits(1) => 
        \sa[13]\, rowbits(0) => VCC_net_1, sa(13) => nc2, sa(12)
         => nc1, sa(11) => sa(11), sa(10) => sa(10), sa(9) => 
        sa(9), sa(8) => sa(8), sa(7) => sa(7), sa(6) => sa(6), 
        sa(5) => sa(5), sa(4) => sa(4), sa(3) => sa(3), sa(2) => 
        sa(2), sa(1) => sa(1), sa(0) => sa(0), ba(1) => ba(1), 
        ba(0) => ba(0), cs_n(0) => cs_n(0), clk => clk, reset_n
         => reset_n, sd_init => \sa[13]\, r_req => \r_req_i\, 
        w_req => \w_req_i\, auto_pch => \sa[13]\, rf_req => 
        \rf_req\, p_req => p_req, m_req => \m_req\, 
        m_req_dll_reset => \sa[13]\, em_req => \sa[13]\, cl_half
         => \sa[13]\, regdimm => \sa[13]\, dqm_wr_bterm => 
        dqm_wr_bterm, rw_ack => rw_ack, s_ack => s_ack, r_valid
         => r_valid, w_valid => w_valid, d_req => OPEN, oe => oe, 
        cke => cke, ras_n => ras_n, cas_n => cas_n, we_n => we_n);
    
    \m_shift[8]\ : SLE
      port map(D => \m_shift[9]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => p_req);
    
    \timer[13]\ : SLE
      port map(D => \timer_p.timer_6[13]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[13]_net_1\);
    
    \init.un5_timer_reset\ : CFG3
      generic map(INIT => x"EC")

      port map(A => s_ack, B => \timer_reset\, C => 
        \start_delay_done\, Y => \init.un5_timer_reset_net_1\);
    
    \timer_p.timer_reset_2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \timer_p.timer_reset_2_9_net_1\, B => 
        \timer_p.timer_reset_2_12_net_1\, C => 
        \timer_p.timer_reset_2_11_net_1\, D => 
        \timer_p.timer_reset_2_10_net_1\, Y => 
        \timer_p.timer_reset_2_net_1\);
    
    \timer[14]\ : SLE
      port map(D => \timer_p.timer_6[14]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[14]_net_1\);
    
    un4_timer_cry_7 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[7]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_6\, S => 
        un4_timer_cry_7_S, Y => OPEN, FCO => \un4_timer_cry_7\);
    
    \timer_RNO[14]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_14_S, Y => \timer_p.timer_6[14]\);
    
    \timer[7]\ : SLE
      port map(D => \timer_p.timer_6[7]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[7]_net_1\);
    
    \timer[10]\ : SLE
      port map(D => \timer_p.timer_6[10]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[10]_net_1\);
    
    \r_shift[1]\ : SLE
      port map(D => \r_shift[2]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[1]_net_1\);
    
    \timer[5]\ : SLE
      port map(D => \timer_p.timer_6[5]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[5]_net_1\);
    
    \timer_RNO[8]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_8_S, Y => \timer_p.timer_6[8]\);
    
    rf_req : SLE
      port map(D => \r_shift[0]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \rf_req\);
    
    \timer_RNO[3]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_3_S, Y => \timer_p.timer_6[3]\);
    
    \timer[12]\ : SLE
      port map(D => \timer_p.timer_6[12]\, CLK => clk, EN => 
        VCC_net_1, ALn => reset_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => \sa[13]\, LAT => \sa[13]\, Q => 
        \timer[12]_net_1\);
    
    \r_shift[6]\ : SLE
      port map(D => \r_shift[7]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[6]_net_1\);
    
    \m_shift[6]\ : SLE
      port map(D => \m_shift[7]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[6]_net_1\);
    
    \r_shift[0]\ : SLE
      port map(D => \r_shift[1]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[0]_net_1\);
    
    \r_shift[4]\ : SLE
      port map(D => \r_shift[5]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[4]_net_1\);
    
    \r_shift[5]\ : SLE
      port map(D => \r_shift[6]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[5]_net_1\);
    
    un4_timer_cry_2 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[2]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_1\, S => 
        un4_timer_cry_2_S, Y => OPEN, FCO => \un4_timer_cry_2\);
    
    inited_RNO : CFG2
      generic map(INIT => x"E")

      port map(A => \dqm_init_p.un6_m_req_net_1\, B => \load\, Y
         => un1_dll_holdoff_en2_i);
    
    un4_timer_cry_3 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[3]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_2\, S => 
        un4_timer_cry_3_S, Y => OPEN, FCO => \un4_timer_cry_3\);
    
    \timer_p.timer_reset_2_12\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \load\, B => \timer_p.timer_reset_2_0_net_1\, 
        C => \timer[14]_net_1\, D => \timer[0]_net_1\, Y => 
        \timer_p.timer_reset_2_12_net_1\);
    
    r_req_i : CFG2
      generic map(INIT => x"8")

      port map(A => r_req, B => \inited\, Y => \r_req_i\);
    
    \timer_p.timer_reset_2_9\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \timer[5]_net_1\, B => \timer[4]_net_1\, C
         => \timer[3]_net_1\, D => \timer[2]_net_1\, Y => 
        \timer_p.timer_reset_2_9_net_1\);
    
    dqm_init : SLE
      port map(D => \sa[13]\, CLK => clk, EN => 
        \dqm_init_p.un6_m_req_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \dqm_init\);
    
    \timer_RNO[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_2_S, Y => \timer_p.timer_6[2]\);
    
    \m_shift[1]\ : SLE
      port map(D => \m_shift[2]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[1]_net_1\);
    
    un4_timer_s_15 : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \timer[15]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_14\, S => 
        un4_timer_s_15_S, Y => OPEN, FCO => OPEN);
    
    \m_shift[4]\ : SLE
      port map(D => \m_shift[5]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \m_shift[4]_net_1\);
    
    dqm_init_d0 : SLE
      port map(D => \dqm_init\, CLK => clk, EN => VCC_net_1, ALn
         => reset_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \sa[13]\, LAT => \sa[13]\, Q => \dqm_init_d0\);
    
    \r_shift_0[9]\ : CFG4
      generic map(INIT => x"0F78")

      port map(A => \start_delay_done\, B => s_ack, C => 
        \r_shift[9]_net_1\, D => \timer_reset\, Y => 
        \r_shift_0[9]_net_1\);
    
    un4_timer_cry_12 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[12]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_11\, S => 
        un4_timer_cry_12_S, Y => OPEN, FCO => \un4_timer_cry_12\);
    
    \timer_p.timer_6_f0[7]\ : CFG3
      generic map(INIT => x"32")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_7_S, Y => \timer_p.timer_6[7]\);
    
    un4_timer_cry_11 : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \timer[11]_net_1\, C => 
        \sa[13]\, D => \sa[13]\, FCI => \un4_timer_cry_10\, S => 
        un4_timer_cry_11_S, Y => OPEN, FCO => \un4_timer_cry_11\);
    
    w_req_i : CFG2
      generic map(INIT => x"8")

      port map(A => w_req, B => \inited\, Y => \w_req_i\);
    
    \timer_p.timer_6_f0[4]\ : CFG3
      generic map(INIT => x"32")

      port map(A => \load\, B => \timer_reset\, C => 
        un4_timer_cry_4_S, Y => \timer_p.timer_6[4]\);
    
    \r_shift[7]\ : SLE
      port map(D => \r_shift[8]_net_1\, CLK => clk, EN => 
        \init.un5_timer_reset_net_1\, ALn => reset_n, ADn => 
        \sa[13]\, SLn => VCC_net_1, SD => \sa[13]\, LAT => 
        \sa[13]\, Q => \r_shift[7]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CORESDR is

    port( RADDR    : in    std_logic_vector(30 downto 0);
          B_SIZE   : in    std_logic_vector(3 downto 0);
          RAS      : in    std_logic_vector(3 downto 0);
          RCD      : in    std_logic_vector(2 downto 0);
          RRD      : in    std_logic_vector(1 downto 0);
          RP       : in    std_logic_vector(2 downto 0);
          RC       : in    std_logic_vector(3 downto 0);
          RFC      : in    std_logic_vector(3 downto 0);
          WR       : in    std_logic_vector(1 downto 0);
          MRD      : in    std_logic_vector(2 downto 0);
          CL       : in    std_logic_vector(2 downto 0);
          BL       : in    std_logic_vector(1 downto 0);
          DELAY    : in    std_logic_vector(15 downto 0);
          REF      : in    std_logic_vector(15 downto 0);
          COLBITS  : in    std_logic_vector(2 downto 0);
          ROWBITS  : in    std_logic_vector(1 downto 0);
          SA       : out   std_logic_vector(13 downto 0);
          BA       : out   std_logic_vector(1 downto 0);
          CS_N     : out   std_logic_vector(0 to 0);
          CLK      : in    std_logic;
          RESET_N  : in    std_logic;
          R_REQ    : in    std_logic;
          W_REQ    : in    std_logic;
          AUTO_PCH : in    std_logic;
          SD_INIT  : in    std_logic;
          REGDIMM  : in    std_logic;
          RW_ACK   : out   std_logic;
          R_VALID  : out   std_logic;
          D_REQ    : out   std_logic;
          W_VALID  : out   std_logic;
          OE       : out   std_logic;
          DQM      : out   std_logic;
          CKE      : out   std_logic;
          RAS_N    : out   std_logic;
          CAS_N    : out   std_logic;
          WE_N     : out   std_logic
        );

end CORESDR;

architecture DEF_ARCH of CORESDR is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component fastinit
    port( raddr    : in    std_logic_vector(30 downto 0) := (others => 'U');
          b_size   : in    std_logic_vector(3 downto 0) := (others => 'U');
          ras      : in    std_logic_vector(3 downto 0) := (others => 'U');
          rcd      : in    std_logic_vector(2 downto 0) := (others => 'U');
          rrd      : in    std_logic_vector(1 downto 0) := (others => 'U');
          rp       : in    std_logic_vector(2 downto 0) := (others => 'U');
          rc       : in    std_logic_vector(3 downto 0) := (others => 'U');
          rfc      : in    std_logic_vector(3 downto 0) := (others => 'U');
          wr       : in    std_logic_vector(1 downto 0) := (others => 'U');
          mrd      : in    std_logic_vector(2 downto 0) := (others => 'U');
          cl       : in    std_logic_vector(2 downto 0) := (others => 'U');
          bl       : in    std_logic_vector(1 downto 0) := (others => 'U');
          ds       : in    std_logic_vector(1 downto 0) := (others => 'U');
          delay    : in    std_logic_vector(15 downto 0) := (others => 'U');
          ref      : in    std_logic_vector(15 downto 0) := (others => 'U');
          colbits  : in    std_logic_vector(2 downto 0) := (others => 'U');
          rowbits  : in    std_logic_vector(1 downto 0) := (others => 'U');
          sa       : out   std_logic_vector(13 downto 0);
          ba       : out   std_logic_vector(1 downto 0);
          cs_n     : out   std_logic_vector(0 to 0);
          clk      : in    std_logic := 'U';
          reset_n  : in    std_logic := 'U';
          r_req    : in    std_logic := 'U';
          w_req    : in    std_logic := 'U';
          auto_pch : in    std_logic := 'U';
          sd_init  : in    std_logic := 'U';
          cl_half  : in    std_logic := 'U';
          regdimm  : in    std_logic := 'U';
          rw_ack   : out   std_logic;
          r_valid  : out   std_logic;
          d_req    : out   std_logic;
          w_valid  : out   std_logic;
          oe       : out   std_logic;
          dqm      : out   std_logic;
          cke      : out   std_logic;
          ras_n    : out   std_logic;
          cas_n    : out   std_logic;
          we_n     : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \r_req_in\, \w_req_in\, \SA[13]\, rw_ack_i, r_valid_i, 
        w_valid_i, \sa_i[0]\, \sa_i[1]\, \sa_i[2]\, \sa_i[3]\, 
        \sa_i[4]\, \sa_i[5]\, \sa_i[6]\, \sa_i[7]\, \sa_i[8]\, 
        \sa_i[9]\, \sa_i[10]\, \sa_i[11]\, \ba_i[0]\, \ba_i[1]\, 
        \cs_n_i[0]\, dqm_i, cke_i, ras_n_i, cas_n_i, we_n_i, 
        VCC_net_1, \r_req_i\, \w_req_i\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : fastinit
	Use entity work.fastinit(DEF_ARCH);
begin 

    SA(13) <= \SA[13]\;
    SA(12) <= \SA[13]\;
    D_REQ <= \SA[13]\;

    \BA[1]\ : SLE
      port map(D => \ba_i[1]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => BA(1));
    
    \WE_N\ : SLE
      port map(D => we_n_i, CLK => CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => WE_N);
    
    \SA[7]\ : SLE
      port map(D => \sa_i[7]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(7));
    
    \CS_N[0]\ : SLE
      port map(D => \cs_n_i[0]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => CS_N(0));
    
    \RW_ACK\ : SLE
      port map(D => rw_ack_i, CLK => CLK, EN => VCC_net_1, ALn
         => RESET_N, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => RW_ACK);
    
    w_req_in : CFG2
      generic map(INIT => x"8")

      port map(A => W_REQ, B => \w_req_i\, Y => \w_req_in\);
    
    \GND\ : GND
      port map(Y => \SA[13]\);
    
    \SA[2]\ : SLE
      port map(D => \sa_i[2]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(2));
    
    fastinit_1 : fastinit
      port map(raddr(30) => \SA[13]\, raddr(29) => \SA[13]\, 
        raddr(28) => \SA[13]\, raddr(27) => \SA[13]\, raddr(26)
         => \SA[13]\, raddr(25) => \SA[13]\, raddr(24) => 
        \SA[13]\, raddr(23) => \SA[13]\, raddr(22) => RADDR(22), 
        raddr(21) => RADDR(21), raddr(20) => RADDR(20), raddr(19)
         => RADDR(19), raddr(18) => RADDR(18), raddr(17) => 
        RADDR(17), raddr(16) => RADDR(16), raddr(15) => RADDR(15), 
        raddr(14) => RADDR(14), raddr(13) => RADDR(13), raddr(12)
         => RADDR(12), raddr(11) => RADDR(11), raddr(10) => 
        RADDR(10), raddr(9) => RADDR(9), raddr(8) => RADDR(8), 
        raddr(7) => RADDR(7), raddr(6) => RADDR(6), raddr(5) => 
        RADDR(5), raddr(4) => RADDR(4), raddr(3) => RADDR(3), 
        raddr(2) => RADDR(2), raddr(1) => RADDR(1), raddr(0) => 
        RADDR(0), b_size(3) => \SA[13]\, b_size(2) => B_SIZE(2), 
        b_size(1) => B_SIZE(1), b_size(0) => B_SIZE(0), ras(3)
         => \SA[13]\, ras(2) => \SA[13]\, ras(1) => VCC_net_1, 
        ras(0) => \SA[13]\, rcd(2) => \SA[13]\, rcd(1) => 
        VCC_net_1, rcd(0) => \SA[13]\, rrd(1) => VCC_net_1, 
        rrd(0) => \SA[13]\, rp(2) => \SA[13]\, rp(1) => VCC_net_1, 
        rp(0) => VCC_net_1, rc(3) => VCC_net_1, rc(2) => \SA[13]\, 
        rc(1) => \SA[13]\, rc(0) => \SA[13]\, rfc(3) => VCC_net_1, 
        rfc(2) => \SA[13]\, rfc(1) => \SA[13]\, rfc(0) => 
        VCC_net_1, wr(1) => VCC_net_1, wr(0) => \SA[13]\, mrd(2)
         => \SA[13]\, mrd(1) => VCC_net_1, mrd(0) => \SA[13]\, 
        cl(2) => \SA[13]\, cl(1) => VCC_net_1, cl(0) => \SA[13]\, 
        bl(1) => VCC_net_1, bl(0) => VCC_net_1, ds(1) => \SA[13]\, 
        ds(0) => \SA[13]\, delay(15) => \SA[13]\, delay(14) => 
        \SA[13]\, delay(13) => \SA[13]\, delay(12) => VCC_net_1, 
        delay(11) => VCC_net_1, delay(10) => \SA[13]\, delay(9)
         => VCC_net_1, delay(8) => \SA[13]\, delay(7) => 
        VCC_net_1, delay(6) => \SA[13]\, delay(5) => \SA[13]\, 
        delay(4) => VCC_net_1, delay(3) => \SA[13]\, delay(2) => 
        \SA[13]\, delay(1) => \SA[13]\, delay(0) => \SA[13]\, 
        ref(15) => \SA[13]\, ref(14) => \SA[13]\, ref(13) => 
        \SA[13]\, ref(12) => VCC_net_1, ref(11) => \SA[13]\, 
        ref(10) => \SA[13]\, ref(9) => \SA[13]\, ref(8) => 
        \SA[13]\, ref(7) => \SA[13]\, ref(6) => \SA[13]\, ref(5)
         => \SA[13]\, ref(4) => \SA[13]\, ref(3) => \SA[13]\, 
        ref(2) => \SA[13]\, ref(1) => \SA[13]\, ref(0) => 
        \SA[13]\, colbits(2) => \SA[13]\, colbits(1) => VCC_net_1, 
        colbits(0) => VCC_net_1, rowbits(1) => \SA[13]\, 
        rowbits(0) => VCC_net_1, sa(13) => nc2, sa(12) => nc1, 
        sa(11) => \sa_i[11]\, sa(10) => \sa_i[10]\, sa(9) => 
        \sa_i[9]\, sa(8) => \sa_i[8]\, sa(7) => \sa_i[7]\, sa(6)
         => \sa_i[6]\, sa(5) => \sa_i[5]\, sa(4) => \sa_i[4]\, 
        sa(3) => \sa_i[3]\, sa(2) => \sa_i[2]\, sa(1) => 
        \sa_i[1]\, sa(0) => \sa_i[0]\, ba(1) => \ba_i[1]\, ba(0)
         => \ba_i[0]\, cs_n(0) => \cs_n_i[0]\, clk => CLK, 
        reset_n => RESET_N, r_req => \r_req_in\, w_req => 
        \w_req_in\, auto_pch => \SA[13]\, sd_init => \SA[13]\, 
        cl_half => \SA[13]\, regdimm => \SA[13]\, rw_ack => 
        rw_ack_i, r_valid => r_valid_i, d_req => OPEN, w_valid
         => w_valid_i, oe => OE, dqm => dqm_i, cke => cke_i, 
        ras_n => ras_n_i, cas_n => cas_n_i, we_n => we_n_i);
    
    \CAS_N\ : SLE
      port map(D => cas_n_i, CLK => CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => CAS_N);
    
    w_req_i : SLE
      port map(D => W_REQ, CLK => CLK, EN => VCC_net_1, ALn => 
        RESET_N, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => \w_req_i\);
    
    \SA[0]\ : SLE
      port map(D => \sa_i[0]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(0));
    
    \W_VALID\ : SLE
      port map(D => w_valid_i, CLK => CLK, EN => VCC_net_1, ALn
         => RESET_N, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => W_VALID);
    
    \SA[3]\ : SLE
      port map(D => \sa_i[3]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(3));
    
    \SA[6]\ : SLE
      port map(D => \sa_i[6]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(6));
    
    \R_VALID\ : SLE
      port map(D => r_valid_i, CLK => CLK, EN => VCC_net_1, ALn
         => RESET_N, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => R_VALID);
    
    \RAS_N\ : SLE
      port map(D => ras_n_i, CLK => CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => RAS_N);
    
    \SA[10]\ : SLE
      port map(D => \sa_i[10]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(10));
    
    \DQM\ : SLE
      port map(D => dqm_i, CLK => CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => DQM);
    
    \SA[4]\ : SLE
      port map(D => \sa_i[4]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(4));
    
    \BA[0]\ : SLE
      port map(D => \ba_i[0]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => BA(0));
    
    \SA[5]\ : SLE
      port map(D => \sa_i[5]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(5));
    
    \SA[1]\ : SLE
      port map(D => \sa_i[1]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(1));
    
    r_req_in : CFG2
      generic map(INIT => x"8")

      port map(A => R_REQ, B => \r_req_i\, Y => \r_req_in\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \CKE\ : SLE
      port map(D => cke_i, CLK => CLK, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => CKE);
    
    \SA[11]\ : SLE
      port map(D => \sa_i[11]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(11));
    
    r_req_i : SLE
      port map(D => R_REQ, CLK => CLK, EN => VCC_net_1, ALn => 
        RESET_N, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => \r_req_i\);
    
    \SA[8]\ : SLE
      port map(D => \sa_i[8]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(8));
    
    \SA[9]\ : SLE
      port map(D => \sa_i[9]\, CLK => CLK, EN => VCC_net_1, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        \SA[13]\, LAT => \SA[13]\, Q => SA(9));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CORESDR_AXI is

    port( COREAXI_0_AXImslave16_AWSIZE       : in    std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_ARSIZE       : in    std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_WDATA        : in    std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_AWADDR       : in    std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_ARADDR       : in    std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_WSTRB        : in    std_logic_vector(7 downto 0);
          DQM_c                              : out   std_logic_vector(1 downto 0);
          sdr_datain_reg                     : out   std_logic_vector(15 downto 0);
          SA_c                               : out   std_logic_vector(11 downto 0);
          BA_c                               : out   std_logic_vector(1 downto 0);
          DQ_in                              : in    std_logic_vector(15 downto 0);
          COREAXI_0_AXImslave16_RDATA_m_8    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58   : out   std_logic;
          COREAXI_0_AXImslave16_ARBURST_0    : in    std_logic;
          CS_N_c_0                           : out   std_logic;
          axi_state_0                        : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_0      : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_3      : out   std_logic;
          RDATA_reg_0                        : out   std_logic;
          RDATA_reg_3                        : out   std_logic;
          N_8_i                              : out   std_logic;
          N_23                               : in    std_logic;
          N_3169_i                           : out   std_logic;
          N_77_mux_i                         : out   std_logic;
          N_76_mux_i                         : out   std_logic;
          N_75_mux_i                         : out   std_logic;
          N_69_mux_i                         : out   std_logic;
          N_68_mux_i                         : out   std_logic;
          N_67_mux_i                         : out   std_logic;
          N_72_mux_i                         : out   std_logic;
          N_71_mux_i                         : out   std_logic;
          N_70_mux_i                         : out   std_logic;
          N_80_mux_i                         : out   std_logic;
          N_79_mux_i                         : out   std_logic;
          N_78_mux_i                         : out   std_logic;
          N_3297                             : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID : in    std_logic;
          N_3170_i                           : out   std_logic;
          COREAXI_0_AXImslave16_AWVALID      : in    std_logic;
          N_39                               : out   std_logic;
          WREADY_SI16_i                      : out   std_logic;
          COREAXI_0_AXImslave16_WVALID       : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID      : in    std_logic;
          i22_mux_2_i                        : out   std_logic;
          i22_mux_3_i                        : out   std_logic;
          i22_mux_4_i                        : out   std_logic;
          i22_mux_5_i                        : out   std_logic;
          i17_mux_2_i                        : out   std_logic;
          i17_mux_i                          : out   std_logic;
          i17_mux_0_i                        : out   std_logic;
          i17_mux_1_i                        : out   std_logic;
          i22_mux_i                          : out   std_logic;
          i22_mux_0_i                        : out   std_logic;
          i22_mux_1_i                        : out   std_logic;
          N_389                              : out   std_logic;
          N_3064_i                           : out   std_logic;
          N_3066_i                           : out   std_logic;
          N_3092_i                           : out   std_logic;
          N_3094_i                           : out   std_logic;
          N_3096_i                           : out   std_logic;
          N_3098_i                           : out   std_logic;
          N_3100_i                           : out   std_logic;
          N_3102_i                           : out   std_logic;
          N_74                               : out   std_logic;
          N_3167_i                           : in    std_logic;
          WE_N_c                             : out   std_logic;
          RAS_N_c                            : out   std_logic;
          un1_top_sb_0_3_i_i                 : out   std_logic;
          CKE_c                              : out   std_logic;
          CAS_N_c                            : out   std_logic;
          COREAXI_0_AXImslave16_BVALID       : out   std_logic;
          COREAXI_0_AXImslave16_AWREADY      : out   std_logic;
          COREAXI_0_AXImslave16_ARREADY      : out   std_logic;
          WREADY_SI16                        : out   std_logic;
          SDRCLK_c                           : in    std_logic;
          MSS_READY                          : in    std_logic
        );

end CORESDR_AXI;

architecture DEF_ARCH of CORESDR_AXI is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CORESDR
    port( RADDR    : in    std_logic_vector(30 downto 0) := (others => 'U');
          B_SIZE   : in    std_logic_vector(3 downto 0) := (others => 'U');
          RAS      : in    std_logic_vector(3 downto 0) := (others => 'U');
          RCD      : in    std_logic_vector(2 downto 0) := (others => 'U');
          RRD      : in    std_logic_vector(1 downto 0) := (others => 'U');
          RP       : in    std_logic_vector(2 downto 0) := (others => 'U');
          RC       : in    std_logic_vector(3 downto 0) := (others => 'U');
          RFC      : in    std_logic_vector(3 downto 0) := (others => 'U');
          WR       : in    std_logic_vector(1 downto 0) := (others => 'U');
          MRD      : in    std_logic_vector(2 downto 0) := (others => 'U');
          CL       : in    std_logic_vector(2 downto 0) := (others => 'U');
          BL       : in    std_logic_vector(1 downto 0) := (others => 'U');
          DELAY    : in    std_logic_vector(15 downto 0) := (others => 'U');
          REF      : in    std_logic_vector(15 downto 0) := (others => 'U');
          COLBITS  : in    std_logic_vector(2 downto 0) := (others => 'U');
          ROWBITS  : in    std_logic_vector(1 downto 0) := (others => 'U');
          SA       : out   std_logic_vector(13 downto 0);
          BA       : out   std_logic_vector(1 downto 0);
          CS_N     : out   std_logic_vector(0 to 0);
          CLK      : in    std_logic := 'U';
          RESET_N  : in    std_logic := 'U';
          R_REQ    : in    std_logic := 'U';
          W_REQ    : in    std_logic := 'U';
          AUTO_PCH : in    std_logic := 'U';
          SD_INIT  : in    std_logic := 'U';
          REGDIMM  : in    std_logic := 'U';
          RW_ACK   : out   std_logic;
          R_VALID  : out   std_logic;
          D_REQ    : out   std_logic;
          W_VALID  : out   std_logic;
          OE       : out   std_logic;
          DQM      : out   std_logic;
          CKE      : out   std_logic;
          RAS_N    : out   std_logic;
          CAS_N    : out   std_logic;
          WE_N     : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sdr_dataout_reg[14]_net_1\, VCC_net_1, GND_net_1, 
        \sdr_dataout_reg[15]_net_1\, \sdr_dataout_reg[0]_net_1\, 
        \sdr_dataout_reg[1]_net_1\, \sdr_dataout_reg[2]_net_1\, 
        \sdr_dataout_reg[3]_net_1\, \sdr_dataout_reg[4]_net_1\, 
        \sdr_dataout_reg[5]_net_1\, \sdr_dataout_reg[6]_net_1\, 
        \sdr_dataout_reg[7]_net_1\, \sdr_dataout_reg[8]_net_1\, 
        \sdr_dataout_reg[9]_net_1\, \sdr_dataout_reg[10]_net_1\, 
        \sdr_dataout_reg[11]_net_1\, \sdr_dataout_reg[12]_net_1\, 
        \sdr_dataout_reg[13]_net_1\, \SA_i[2]\, \SA_i[3]\, 
        \SA_i[4]\, \SA_i[5]\, \SA_i[6]\, \SA_i[7]\, \SA_i[8]\, 
        \SA_i[9]\, \SA_i[10]\, \SA_i[11]\, \sdr_datain[5]\, 
        \sdr_datain[6]\, \sdr_datain[7]\, \sdr_datain[8]\, 
        \sdr_datain[9]\, \sdr_datain[10]\, \sdr_datain[11]\, 
        \sdr_datain[12]\, \sdr_datain[13]\, \sdr_datain[14]\, 
        \sdr_datain[15]\, \BA_i[0]\, \BA_i[1]\, \SA_i[0]\, 
        \SA_i[1]\, \sdr_count[2]_net_1\, N_3278_i, 
        \sdr_count[3]_net_1\, N_3277_i, \axi_count[0]_net_1\, 
        N_3276_i, \axi_count[1]_net_1\, N_3273_i, 
        \axi_count[2]_net_1\, N_3272_i, \axi_count[3]_net_1\, 
        N_3271_i, \sdr_datain[0]\, \sdr_datain[1]\, 
        \sdr_datain[2]\, \sdr_datain[3]\, \sdr_datain[4]\, 
        \raddr_reg[18]_net_1\, \raddr_reg_9[18]_net_1\, 
        \raddr_reg[19]_net_1\, \raddr_reg_9[19]_net_1\, 
        \raddr_reg[20]_net_1\, \raddr_reg_9[20]_net_1\, 
        \raddr_reg[21]_net_1\, \raddr_reg_9[21]_net_1\, 
        \raddr_reg[22]_net_1\, \raddr_reg_9[22]_net_1\, 
        \sdr_count[0]_net_1\, N_3280_i, \sdr_count[1]_net_1\, 
        N_3279_i, \raddr_reg[3]_net_1\, \raddr_reg_9[3]_net_1\, 
        \raddr_reg[4]_net_1\, \raddr_reg_9[4]_net_1\, 
        \raddr_reg[5]_net_1\, \raddr_reg_9[5]_net_1\, 
        \raddr_reg[6]_net_1\, \raddr_reg_9[6]_net_1\, 
        \raddr_reg[7]_net_1\, \raddr_reg_9[7]_net_1\, 
        \raddr_reg[8]_net_1\, \raddr_reg_9[8]_net_1\, 
        \raddr_reg[9]_net_1\, \raddr_reg_9[9]_net_1\, 
        \raddr_reg[10]_net_1\, \raddr_reg_9[10]_net_1\, 
        \raddr_reg[11]_net_1\, \raddr_reg_9[11]_net_1\, 
        \raddr_reg[12]_net_1\, \raddr_reg_9[12]_net_1\, 
        \raddr_reg[13]_net_1\, \raddr_reg_9[13]_net_1\, 
        \raddr_reg[14]_net_1\, \raddr_reg_9[14]_net_1\, 
        \raddr_reg[15]_net_1\, \raddr_reg_9[15]_net_1\, 
        \raddr_reg[16]_net_1\, \raddr_reg_9[16]_net_1\, 
        \raddr_reg[17]_net_1\, \raddr_reg_9[17]_net_1\, 
        \WSTRB_reg[3]_net_1\, \WREADY_SI16\, \WSTRB_reg[4]_net_1\, 
        \WSTRB_reg[5]_net_1\, \WSTRB_reg[6]_net_1\, 
        \WSTRB_reg[7]_net_1\, \B_SIZE_reg[0]_net_1\, 
        \asize[1]_net_1\, N_295_i, \B_SIZE_reg[1]_net_1\, b_size3, 
        \B_SIZE_reg[2]_net_1\, b_size4, \DQM_i_1[0]_net_1\, 
        \DQM_i_3[1]_net_1\, \raddr_reg[0]_net_1\, 
        \raddr_reg_9[0]_net_1\, \raddr_reg[1]_net_1\, 
        \raddr_reg_9[1]_net_1\, \raddr_reg[2]_net_1\, 
        \raddr_reg_9[2]_net_1\, \RDATA_reg[52]_net_1\, 
        N_190_mux_i, \R_VALID\, \RDATA_reg[53]_net_1\, 
        N_191_mux_i, \RDATA_reg[54]_net_1\, N_192_mux_i, 
        \RDATA_reg[55]_net_1\, N_193_mux_i, \RDATA_reg[56]_net_1\, 
        N_194_mux_i, \RDATA_reg[57]_net_1\, N_195_mux_i, 
        \RDATA_reg[58]_net_1\, N_196_mux_i, \RDATA_reg[59]_net_1\, 
        N_197_mux_i, \RDATA_reg[60]_net_1\, N_198_mux_i, 
        \RDATA_reg[61]_net_1\, N_199_mux_i, \RDATA_reg[62]_net_1\, 
        N_200_mux_i, \RDATA_reg[63]_net_1\, N_201_mux_i, 
        \WSTRB_reg[0]_net_1\, \WSTRB_reg[1]_net_1\, 
        \WSTRB_reg[2]_net_1\, \RDATA_reg[37]_net_1\, 
        \RDATA_regce[32]_net_1\, \RDATA_reg[38]_net_1\, 
        \RDATA_reg[39]_net_1\, \RDATA_reg[40]_net_1\, 
        \RDATA_reg[41]_net_1\, \RDATA_reg[42]_net_1\, 
        \RDATA_reg[44]_net_1\, \RDATA_reg[45]_net_1\, 
        \RDATA_reg[47]_net_1\, \RDATA_reg[48]_net_1\, N_186_mux_i, 
        \RDATA_reg[49]_net_1\, N_187_mux_i, \RDATA_reg[50]_net_1\, 
        N_188_mux_i, \RDATA_reg[51]_net_1\, N_189_mux_i, 
        \RDATA_reg[22]_net_1\, \RDATA_regce[19]_net_1\, 
        \RDATA_reg[23]_net_1\, \RDATA_reg[24]_net_1\, 
        \RDATA_reg[25]_net_1\, \RDATA_reg[26]_net_1\, 
        \RDATA_reg[27]_net_1\, \RDATA_reg[28]_net_1\, 
        \RDATA_reg[29]_net_1\, N_3072_i, \RDATA_reg[30]_net_1\, 
        N_3073_i, \RDATA_reg[31]_net_1\, N_3074_i, 
        \RDATA_reg[32]_net_1\, \RDATA_reg[33]_net_1\, 
        \RDATA_reg[34]_net_1\, \RDATA_reg[35]_net_1\, 
        \RDATA_reg[36]_net_1\, \COREAXI_0_AXImslave16_RDATA[7]\, 
        N_177_mux_i, \COREAXI_0_AXImslave16_RDATA[8]\, 
        N_178_mux_i, \COREAXI_0_AXImslave16_RDATA[9]\, 
        N_179_mux_i, \COREAXI_0_AXImslave16_RDATA[10]\, 
        N_180_mux_i, \COREAXI_0_AXImslave16_RDATA_0\, N_181_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[12]\, N_182_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[13]\, N_183_mux_i, 
        \COREAXI_0_AXImslave16_RDATA_3\, N_184_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[15]\, N_185_mux_i, 
        \RDATA_reg[16]_net_1\, N_3069_i, \RDATA_reg[17]_net_1\, 
        N_3070_i, \RDATA_reg[18]_net_1\, N_3071_i, 
        \RDATA_reg[19]_net_1\, \RDATA_reg[20]_net_1\, 
        \RDATA_reg[21]_net_1\, \WDATA_reg[56]_net_1\, 
        \WDATA_mux[56]\, \WDATA_reg[57]_net_1\, \WDATA_mux[57]\, 
        \WDATA_reg[58]_net_1\, \WDATA_mux[58]\, 
        \WDATA_reg[59]_net_1\, \WDATA_mux[59]\, 
        \WDATA_reg[60]_net_1\, \WDATA_mux[60]\, 
        \WDATA_reg[61]_net_1\, \WDATA_mux[61]\, 
        \WDATA_reg[62]_net_1\, \WDATA_mux[62]\, 
        \WDATA_reg[63]_net_1\, \WDATA_mux[63]\, 
        \COREAXI_0_AXImslave16_RDATA[0]\, N_170_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[1]\, N_171_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[2]\, N_172_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[3]\, N_173_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[4]\, N_174_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[5]\, N_175_mux_i, 
        \COREAXI_0_AXImslave16_RDATA[6]\, N_176_mux_i, 
        \WDATA_reg[41]_net_1\, \WDATA_mux[41]\, 
        \WDATA_reg[42]_net_1\, \WDATA_mux[42]\, 
        \WDATA_reg[43]_net_1\, \WDATA_mux[43]\, 
        \WDATA_reg[44]_net_1\, \WDATA_mux[44]\, 
        \WDATA_reg[45]_net_1\, \WDATA_mux[45]\, 
        \WDATA_reg[46]_net_1\, \WDATA_mux[46]\, 
        \WDATA_reg[47]_net_1\, \WDATA_mux[47]\, 
        \WDATA_reg[48]_net_1\, \WDATA_mux[48]\, 
        \WDATA_reg[49]_net_1\, \WDATA_mux[49]\, 
        \WDATA_reg[50]_net_1\, \WDATA_mux[50]\, 
        \WDATA_reg[51]_net_1\, \WDATA_mux[51]\, 
        \WDATA_reg[52]_net_1\, \WDATA_mux[52]\, 
        \WDATA_reg[53]_net_1\, \WDATA_mux[53]\, 
        \WDATA_reg[54]_net_1\, \WDATA_mux[54]\, 
        \WDATA_reg[55]_net_1\, \WDATA_mux[55]\, 
        \WDATA_reg[26]_net_1\, \WDATA_mux[26]\, 
        \WDATA_reg[27]_net_1\, \WDATA_mux[27]\, 
        \WDATA_reg[28]_net_1\, \WDATA_mux[28]\, 
        \WDATA_reg[29]_net_1\, \WDATA_mux[29]\, 
        \WDATA_reg[30]_net_1\, \WDATA_mux[30]\, 
        \WDATA_reg[31]_net_1\, \WDATA_mux[31]\, 
        \WDATA_reg[32]_net_1\, \WDATA_mux[32]\, 
        \WDATA_reg[33]_net_1\, \WDATA_mux[33]\, 
        \WDATA_reg[34]_net_1\, \WDATA_mux[34]\, 
        \WDATA_reg[35]_net_1\, \WDATA_mux[35]\, 
        \WDATA_reg[36]_net_1\, \WDATA_mux[36]\, 
        \WDATA_reg[37]_net_1\, \WDATA_mux[37]\, 
        \WDATA_reg[38]_net_1\, \WDATA_mux[38]\, 
        \WDATA_reg[39]_net_1\, \WDATA_mux[39]\, 
        \WDATA_reg[40]_net_1\, \WDATA_mux[40]\, 
        \WDATA_reg[11]_net_1\, \WDATA_mux[11]\, 
        \WDATA_reg[12]_net_1\, \WDATA_mux[12]\, 
        \WDATA_reg[13]_net_1\, \WDATA_mux[13]\, 
        \WDATA_reg[14]_net_1\, \WDATA_mux[14]\, 
        \WDATA_reg[15]_net_1\, \WDATA_mux[15]\, 
        \WDATA_reg[16]_net_1\, \WDATA_mux[16]\, 
        \WDATA_reg[17]_net_1\, \WDATA_mux[17]\, 
        \WDATA_reg[18]_net_1\, \WDATA_mux[18]\, 
        \WDATA_reg[19]_net_1\, \WDATA_mux[19]\, 
        \WDATA_reg[20]_net_1\, \WDATA_mux[20]\, 
        \WDATA_reg[21]_net_1\, \WDATA_mux[21]\, 
        \WDATA_reg[22]_net_1\, \WDATA_mux[22]\, 
        \WDATA_reg[23]_net_1\, \WDATA_mux[23]\, 
        \WDATA_reg[24]_net_1\, \WDATA_mux[24]\, 
        \WDATA_reg[25]_net_1\, \WDATA_mux[25]\, 
        \asize_reg[0]_net_1\, \asize_reg_134\, 
        \asize_reg[1]_net_1\, \asize_reg_135\, 
        \WDATA_reg[0]_net_1\, \WDATA_mux[0]\, 
        \WDATA_reg[1]_net_1\, \WDATA_mux[1]\, 
        \WDATA_reg[2]_net_1\, \WDATA_mux[2]\, 
        \WDATA_reg[3]_net_1\, \WDATA_mux[3]\, 
        \WDATA_reg[4]_net_1\, \WDATA_mux[4]\, 
        \WDATA_reg[5]_net_1\, \WDATA_mux[5]\, 
        \WDATA_reg[6]_net_1\, \WDATA_mux[6]\, 
        \WDATA_reg[7]_net_1\, \WDATA_mux[7]\, 
        \WDATA_reg[8]_net_1\, \WDATA_mux[8]\, 
        \WDATA_reg[9]_net_1\, \WDATA_mux[9]\, 
        \WDATA_reg[10]_net_1\, \WDATA_mux[10]\, \R_VALID_reg\, 
        R_VALID_i, \axi_state[0]_net_1\, \axi_state_ns[9]_net_1\, 
        \axi_state[9]_net_1\, \axi_state_ns[0]\, 
        \COREAXI_0_AXImslave16_ARREADY\, \axi_state_ns[1]_net_1\, 
        \COREAXI_0_AXImslave16_AWREADY\, \axi_state_ns[2]_net_1\, 
        \axi_state_0\, \axi_state_ns[3]_net_1\, 
        \axi_state[5]_net_1\, N_308_i, 
        \COREAXI_0_AXImslave16_BVALID\, \axi_state_ns[5]\, 
        \axi_state[3]_net_1\, N_311_i, \axi_state[2]_net_1\, 
        \axi_state_ns[7]\, \axi_state[1]_net_1\, 
        \axi_state_ns[8]_net_1\, CAS_N_i, CKE_i, \CS_N_i[0]\, 
        OE_i, RAS_N_i, WE_N_i, raddr_reg_9_2_cry_0, 
        \un1_B_SIZE_reg_0_a2_RNISOQQ1_Y[2]\, 
        \un1_B_SIZE_reg_0_a2[2]_net_1\, N_335_i, 
        \raddr_reg_RNIOTA71[0]_net_1\, raddr_reg_9_2_cry_1, N_750, 
        \un1_B_SIZE_reg_0_a2[1]_net_1\, 
        \raddr_reg_RNIR0B71[1]_net_1\, raddr_reg_9_2_cry_2, N_751, 
        \un1_B_SIZE_reg_0_a2[0]_net_1\, 
        \raddr_reg_RNIU3B71[2]_net_1\, raddr_reg_9_2_cry_3, N_752, 
        \raddr_reg_9_2_axb_3_1\, raddr_reg_9_sn_N_3_i, 
        raddr_reg_9_2_cry_4, N_753, \raddr_reg_9_2_axb_4_1\, 
        raddr_reg_9_2_cry_5, N_754, \raddr_reg_9_2_axb_5_1\, 
        raddr_reg_9_2_cry_6, N_755, \raddr_reg_9_2_axb_6_1\, 
        raddr_reg_9_2_cry_7, N_756, \raddr_reg_9_2_axb_7_1\, 
        raddr_reg_9_2_cry_8, N_757, \raddr_reg_9_2_axb_8_1\, 
        raddr_reg_9_2_cry_9, N_758, \raddr_reg_9_2_axb_9_1\, 
        raddr_reg_9_2_cry_10, N_759, \raddr_reg_9_2_axb_10_1\, 
        raddr_reg_9_2_cry_11, N_760, \raddr_reg_9_2_axb_11_1\, 
        raddr_reg_9_2_cry_12, N_761, \raddr_reg_9_2_axb_12_1\, 
        raddr_reg_9_2_cry_13, N_762, \raddr_reg_9_2_axb_13_1\, 
        raddr_reg_9_2_cry_14, N_763, \raddr_reg_9_2_axb_14_1\, 
        raddr_reg_9_2_cry_15, N_764, \raddr_reg_9_2_axb_15_1\, 
        raddr_reg_9_2_cry_16, N_765, \raddr_reg_9_2_axb_16_1\, 
        raddr_reg_9_2_cry_17, N_766, \raddr_reg_9_2_axb_17_1\, 
        raddr_reg_9_2_cry_18, N_767, \raddr_reg_9_2_axb_18_1\, 
        raddr_reg_9_2_cry_19, N_768, \raddr_reg_9_2_axb_19_1\, 
        raddr_reg_9_2_cry_20, N_769, \raddr_reg_9_2_axb_20_1\, 
        N_771, raddr_reg_9_2_axb_22_1, raddr_reg_9_2_cry_21, 
        N_770, \raddr_reg_9_2_axb_21_1\, N_3281, 
        un1_sdr_count_0_sqmuxa, N_3293, N_3288, WDATA_mux_8_sm0, 
        \WDATA_mux_8_3[7]_net_1\, \WDATA_mux_8_3[6]_net_1\, 
        \WDATA_mux_8_3[5]_net_1\, \WDATA_mux_8_3[4]_net_1\, 
        \WDATA_mux_8_3[3]_net_1\, \WDATA_mux_8_3[2]_net_1\, 
        \WDATA_mux_8_3[1]_net_1\, \WDATA_mux_8_3[0]_net_1\, 
        WDATA_mux_15_sm0, \WDATA_mux_15_3[15]_net_1\, 
        \WDATA_mux_15_3[14]_net_1\, \WDATA_mux_15_3[13]_net_1\, 
        \WDATA_mux_15_3[12]_net_1\, \WDATA_mux_15_3[11]_net_1\, 
        \WDATA_mux_15_3[10]_net_1\, \WDATA_mux_15_3[9]_net_1\, 
        \WDATA_mux_15_3[8]_net_1\, \WDATA_mux_8_m0[0]\, 
        \WDATA_mux_8_0[0]_net_1\, \WDATA_mux_8_0[7]_net_1\, 
        \WDATA_mux_8_0[6]_net_1\, \WDATA_mux_8_0[5]_net_1\, 
        \WDATA_mux_8_0[4]_net_1\, \WDATA_mux_8_0[3]_net_1\, 
        \WDATA_mux_8_0[2]_net_1\, \WDATA_mux_8_0[1]_net_1\, 
        \WDATA_mux_15_0[15]_net_1\, \WDATA_mux_15_0[14]_net_1\, 
        \WDATA_mux_15_0[13]_net_1\, \WDATA_mux_15_0[12]_net_1\, 
        \WDATA_mux_15_0[11]_net_1\, \WDATA_mux_15_0[10]_net_1\, 
        \WDATA_mux_15_0[9]_net_1\, \WDATA_mux_15_0[8]_net_1\, 
        \N_74\, N_3149_2, \N_389\, \raddr_reg_9_2_1_1[1]_net_1\, 
        \COREAXI_0_AXImslave16_RDATA_m_8\, i22_mux_1_i_1_0, 
        i22_mux_1_i_1, \COREAXI_0_AXImslave16_RDATA_m_11\, 
        i22_mux_0_i_1_0, i22_mux_0_i_1, 
        \COREAXI_0_AXImslave16_RDATA_m_12\, i22_mux_i_1_0, 
        i22_mux_i_1, \COREAXI_0_AXImslave16_RDATA_m_13\, 
        i17_mux_1_i_1_0, i17_mux_1_i_1, 
        \COREAXI_0_AXImslave16_RDATA_m_14\, i17_mux_0_i_1_0, 
        i17_mux_0_i_1, \COREAXI_0_AXImslave16_RDATA_m_15\, 
        i17_mux_i_1_0, i17_mux_i_1, 
        \COREAXI_0_AXImslave16_RDATA_m_0\, i17_mux_2_i_1_0, 
        i17_mux_2_i_1, \COREAXI_0_AXImslave16_RDATA_m_4\, 
        i22_mux_5_i_1_0, i22_mux_5_i_1, 
        \COREAXI_0_AXImslave16_RDATA_m_5\, i22_mux_4_i_1_0, 
        i22_mux_4_i_1, \COREAXI_0_AXImslave16_RDATA_m_6\, 
        i22_mux_3_i_1_0, i22_mux_3_i_1, 
        \COREAXI_0_AXImslave16_RDATA_m_7\, i22_mux_2_i_1_0, 
        i22_mux_2_i_1, m30_1_1_2, i58_mux_2, m9_1_1_2, i58_mux, 
        m23_1_2, i58_mux_1, \WSTRB_mux_8_m1_1[0]_net_1\, 
        \un7_wstrb_reg_i_a3\, \WSTRB_mux_8_m1[0]_net_1\, 
        m16_1_1_2, i58_mux_0, \WSTRB_mux_8_m1_1[1]_net_1\, 
        \WSTRB_mux_8_m1[1]_net_1\, \raddr_reg_9_2_1_1[0]_net_1\, 
        \raddr_reg_9_2_1_1[2]_net_1\, \DQM_mux_ns_1_1[1]_net_1\, 
        \WSTRB_mux[3]\, \DQM_mux_ns_1[1]_net_1\, 
        \sdr_count_RNI201B[3]_net_1\, N_3153, N_3144, 
        \DQM_mux[1]\, \DQM_mux_ns_1_1[0]_net_1\, \WSTRB_mux[2]\, 
        \DQM_mux_ns_1[0]_net_1\, N_3154, N_3145, \DQM_mux[0]\, 
        \WDATA_mux_8_1[7]_net_1\, \WDATA_mux_8[7]\, 
        \WDATA_mux_8_1[6]_net_1\, \WDATA_mux_8[6]\, 
        \WDATA_mux_8_1[5]_net_1\, \WDATA_mux_8[5]\, 
        \WDATA_mux_8_1[4]_net_1\, \WDATA_mux_8[4]\, 
        \WDATA_mux_8_1[3]_net_1\, \WDATA_mux_8[3]\, 
        \WDATA_mux_8_1[2]_net_1\, \WDATA_mux_8[2]\, 
        \WDATA_mux_8_1[1]_net_1\, \WDATA_mux_8[1]\, 
        \WDATA_mux_8_1[0]_net_1\, \WDATA_mux_8[0]\, 
        \WDATA_mux_15_1[15]_net_1\, \WDATA_mux_15[15]\, 
        \WDATA_mux_15_1[14]_net_1\, \WDATA_mux_15[14]\, 
        \WDATA_mux_15_1[13]_net_1\, \WDATA_mux_15[13]\, 
        \WDATA_mux_15_1[12]_net_1\, \WDATA_mux_15[12]\, 
        \WDATA_mux_15_1[11]_net_1\, \WDATA_mux_15[11]\, 
        \WDATA_mux_15_1[10]_net_1\, \WDATA_mux_15[10]\, 
        \WDATA_mux_15_1[9]_net_1\, \WDATA_mux_15[9]\, 
        \WDATA_mux_15_1[8]_net_1\, \WDATA_mux_15[8]\, 
        \sdr_datain_3[15]_net_1\, \sdr_datain_1[15]_net_1\, 
        \sdr_datain_2[15]_net_1\, \sdr_datain_0[15]_net_1\, 
        \sdr_datain_3[14]_net_1\, \sdr_datain_1[14]_net_1\, 
        \sdr_datain_2[14]_net_1\, \sdr_datain_0[14]_net_1\, 
        \sdr_datain_3[13]_net_1\, \sdr_datain_1[13]_net_1\, 
        \sdr_datain_2[13]_net_1\, \sdr_datain_0[13]_net_1\, 
        \sdr_datain_3[12]_net_1\, \sdr_datain_1[12]_net_1\, 
        \sdr_datain_2[12]_net_1\, \sdr_datain_0[12]_net_1\, 
        \sdr_datain_3[11]_net_1\, \sdr_datain_1[11]_net_1\, 
        \sdr_datain_2[11]_net_1\, \sdr_datain_0[11]_net_1\, 
        \sdr_datain_3[10]_net_1\, \sdr_datain_1[10]_net_1\, 
        \sdr_datain_2[10]_net_1\, \sdr_datain_0[10]_net_1\, 
        \sdr_datain_3[9]_net_1\, \sdr_datain_1[9]_net_1\, 
        \sdr_datain_2[9]_net_1\, \sdr_datain_0[9]_net_1\, 
        \sdr_datain_3[8]_net_1\, \sdr_datain_1[8]_net_1\, 
        \sdr_datain_2[8]_net_1\, \sdr_datain_0[8]_net_1\, 
        \sdr_datain_3[7]_net_1\, \sdr_datain_1[7]_net_1\, 
        \sdr_datain_2[7]_net_1\, \sdr_datain_0[7]_net_1\, 
        \sdr_datain_3[6]_net_1\, \sdr_datain_1[6]_net_1\, 
        \sdr_datain_2[6]_net_1\, \sdr_datain_0[6]_net_1\, 
        \sdr_datain_3[5]_net_1\, \sdr_datain_1[5]_net_1\, 
        \sdr_datain_2[5]_net_1\, \sdr_datain_0[5]_net_1\, 
        \sdr_datain_3[4]_net_1\, \sdr_datain_1[4]_net_1\, 
        \sdr_datain_2[4]_net_1\, \sdr_datain_0[4]_net_1\, 
        \sdr_datain_3[3]_net_1\, \sdr_datain_1[3]_net_1\, 
        \sdr_datain_2[3]_net_1\, \sdr_datain_0[3]_net_1\, 
        \sdr_datain_3[2]_net_1\, \sdr_datain_1[2]_net_1\, 
        \sdr_datain_2[2]_net_1\, \sdr_datain_0[2]_net_1\, 
        \sdr_datain_3[1]_net_1\, \sdr_datain_1[1]_net_1\, 
        \sdr_datain_2[1]_net_1\, \sdr_datain_0[1]_net_1\, 
        \sdr_datain_3[0]_net_1\, \sdr_datain_1[0]_net_1\, 
        \sdr_datain_2[0]_net_1\, \sdr_datain_0[0]_net_1\, 
        \WSTRB_mux_3_0_a3_0_0[2]_net_1\, 
        \WSTRB_mux_3_0_a3_0_0[3]_net_1\, N_3157, N_3286, N_3141, 
        N_358, W_VALID, N_388, un5_axi_rvalid_i_0, 
        \asize[0]_net_1\, \axi_state_ns_i_0[4]_net_1\, RW_ACK, 
        \axi_state_ns_0_0[7]_net_1\, WSTRB_mux_8_sn_m3_i_a3_1, 
        N_3313, N_3200, N_3326_i, N_3236, N_3207, N_3268, N_3172, 
        N_72, N_343_i, N_3240, \WDATA_mux_31[17]_net_1\, 
        \WDATA_mux_31[18]_net_1\, \WDATA_mux_31[19]_net_1\, 
        \WDATA_mux_31[20]_net_1\, \WDATA_mux_31[21]_net_1\, 
        \WDATA_mux_31[22]_net_1\, \WDATA_mux_31[23]_net_1\, 
        N_3210, \axi_state_ns_0_0[0]_net_1\, 
        \COREAXI_0_AXImslave16_RDATA_m_i_0[51]\, 
        \WDATA_mux_3_0_0[16]_net_1\, un2_sdr_count_NE_0, N_3202, 
        N_71_i, \N_3297\, N_355_i, N_26, 
        \WDATA_mux_3_0_0[5]_net_1\, \WDATA_mux_3_0_0[6]_net_1\, 
        \WDATA_mux_3_0_0[4]_net_1\, \WDATA_mux_3_0_0[7]_net_1\, 
        \WDATA_mux_3_0_0[0]_net_1\, \WDATA_mux_3_0_0[3]_net_1\, 
        \WDATA_mux_3_0_0[1]_net_1\, \WDATA_mux_3_0_0[2]_net_1\, 
        \WDATA_mux_3_0_0[9]_net_1\, \WDATA_mux_3_0_0[8]_net_1\, 
        \WDATA_mux_3_0_0[10]_net_1\, \WDATA_mux_3_0_0[11]_net_1\, 
        \WDATA_mux_3_0_0[12]_net_1\, \WDATA_mux_3_0_0[13]_net_1\, 
        \WDATA_mux_3_0_0[15]_net_1\, \WDATA_mux_3_0_1[14]_net_1\, 
        \un3_r_req_0_0\, N_3299, N_3289, N_338, N_349, N_368, 
        N_3309, dqm_sdr : std_logic;
    signal nc2, nc1 : std_logic;

    for all : CORESDR
	Use entity work.CORESDR(DEF_ARCH);
begin 

    COREAXI_0_AXImslave16_RDATA_m_8 <= 
        \COREAXI_0_AXImslave16_RDATA_m_8\;
    COREAXI_0_AXImslave16_RDATA_m_11 <= 
        \COREAXI_0_AXImslave16_RDATA_m_11\;
    COREAXI_0_AXImslave16_RDATA_m_12 <= 
        \COREAXI_0_AXImslave16_RDATA_m_12\;
    COREAXI_0_AXImslave16_RDATA_m_13 <= 
        \COREAXI_0_AXImslave16_RDATA_m_13\;
    COREAXI_0_AXImslave16_RDATA_m_14 <= 
        \COREAXI_0_AXImslave16_RDATA_m_14\;
    COREAXI_0_AXImslave16_RDATA_m_15 <= 
        \COREAXI_0_AXImslave16_RDATA_m_15\;
    COREAXI_0_AXImslave16_RDATA_m_0 <= 
        \COREAXI_0_AXImslave16_RDATA_m_0\;
    COREAXI_0_AXImslave16_RDATA_m_4 <= 
        \COREAXI_0_AXImslave16_RDATA_m_4\;
    COREAXI_0_AXImslave16_RDATA_m_5 <= 
        \COREAXI_0_AXImslave16_RDATA_m_5\;
    COREAXI_0_AXImslave16_RDATA_m_6 <= 
        \COREAXI_0_AXImslave16_RDATA_m_6\;
    COREAXI_0_AXImslave16_RDATA_m_7 <= 
        \COREAXI_0_AXImslave16_RDATA_m_7\;
    axi_state_0 <= \axi_state_0\;
    COREAXI_0_AXImslave16_RDATA_0 <= 
        \COREAXI_0_AXImslave16_RDATA_0\;
    COREAXI_0_AXImslave16_RDATA_3 <= 
        \COREAXI_0_AXImslave16_RDATA_3\;
    N_3297 <= \N_3297\;
    N_389 <= \N_389\;
    N_74 <= \N_74\;
    COREAXI_0_AXImslave16_BVALID <= 
        \COREAXI_0_AXImslave16_BVALID\;
    COREAXI_0_AXImslave16_AWREADY <= 
        \COREAXI_0_AXImslave16_AWREADY\;
    COREAXI_0_AXImslave16_ARREADY <= 
        \COREAXI_0_AXImslave16_ARREADY\;
    WREADY_SI16 <= \WREADY_SI16\;

    \raddr_reg_RNIU3B71[2]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \raddr_reg[2]_net_1\, B => 
        \raddr_reg_9_2_1_1[2]_net_1\, C => raddr_reg_9_sn_N_3_i, 
        Y => \raddr_reg_RNIU3B71[2]_net_1\);
    
    \axi_count_7_i_o2_0[0]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WVALID, B => 
        \axi_state_0\, C => \axi_state[5]_net_1\, D => N_23, Y
         => N_3281);
    
    \WDATA_reg[34]\ : SLE
      port map(D => \WDATA_mux[34]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[34]_net_1\);
    
    \sdr_datain_0[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[23]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[7]_net_1\);
    
    \sdr_datain_reg[9]\ : SLE
      port map(D => \sdr_datain[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(9));
    
    \DQM_mux_ns[1]\ : CFG4
      generic map(INIT => x"0257")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => N_3153, C
         => N_3144, D => \DQM_mux_ns_1[1]_net_1\, Y => 
        \DQM_mux[1]\);
    
    \sdr_dataout_reg[3]\ : SLE
      port map(D => DQ_in(3), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[3]_net_1\);
    
    \raddr_reg[13]\ : SLE
      port map(D => \raddr_reg_9[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[13]_net_1\);
    
    \WDATA_mux_8_3[3]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(3), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[3]_net_1\);
    
    \axi_state_ns[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \axi_state[2]_net_1\, B => 
        \axi_state[1]_net_1\, C => RW_ACK, D => N_349, Y => 
        \axi_state_ns[8]_net_1\);
    
    \sdr_datain_2[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[8]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[8]_net_1\);
    
    \SA[3]\ : SLE
      port map(D => \SA_i[3]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(3));
    
    \un1_axi_state_4_i_o2[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \axi_state[0]_net_1\, B => 
        \axi_state[1]_net_1\, Y => N_335_i);
    
    \WDATA_mux_8_0[2]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(50), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[2]_net_1\);
    
    un61_axi_state_i_o2 : CFG4
      generic map(INIT => x"FFF7")

      port map(A => N_71_i, B => N_3326_i, C => 
        un2_sdr_count_NE_0, D => N_388, Y => N_343_i);
    
    \WDATA_reg[19]\ : SLE
      port map(D => \WDATA_mux[19]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[19]_net_1\);
    
    \WDATA_mux_3_0_0[16]\ : CFG4
      generic map(INIT => x"80AA")

      port map(A => COREAXI_0_AXImslave16_WDATA(16), B => 
        \asize_reg[1]_net_1\, C => COREAXI_0_AXImslave16_WSTRB(2), 
        D => \N_74\, Y => \WDATA_mux_3_0_0[16]_net_1\);
    
    \sdr_dataout_reg[11]\ : SLE
      port map(D => DQ_in(11), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[11]_net_1\);
    
    \RDATA_reg[4]\ : SLE
      port map(D => N_174_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[4]\);
    
    \WSTRB_mux_8_m1[0]\ : CFG4
      generic map(INIT => x"FAF8")

      port map(A => \WSTRB_mux_8_m1_1[0]_net_1\, B => 
        \un7_wstrb_reg_i_a3\, C => \WSTRB_reg[2]_net_1\, D => 
        \WSTRB_reg[4]_net_1\, Y => \WSTRB_mux_8_m1[0]_net_1\);
    
    \WDATA_mux_3[17]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(17), C => 
        \WDATA_mux_31[17]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[17]\);
    
    \asize_reg_RNIOB215[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_12\, C => i22_mux_i_1_0, D
         => i22_mux_i_1, Y => i22_mux_i);
    
    \WDATA_reg_RNO[37]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(37), 
        Y => \WDATA_mux[37]\);
    
    \sdr_datain_reg_RNO[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[0]_net_1\, C => \sdr_datain_1[0]_net_1\, Y
         => \sdr_datain[0]\);
    
    \raddr_reg[4]\ : SLE
      port map(D => \raddr_reg_9[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[4]_net_1\);
    
    \RDATA_reg_RNIOKCR1[45]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[13]\, B => 
        \RDATA_reg[45]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3064_i);
    
    \un7_1.N_3271_i\ : CFG4
      generic map(INIT => x"00C9")

      port map(A => N_3286, B => \axi_count[3]_net_1\, C => 
        N_3289, D => N_3293, Y => N_3271_i);
    
    \RDATA_reg[63]\ : SLE
      port map(D => N_201_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[63]_net_1\);
    
    \RDATA_reg_RNITOGN1[54]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[54]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_3_i_1);
    
    \sdr_count_9_i_o2[2]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => un1_sdr_count_0_sqmuxa, Y => 
        N_3288);
    
    \RDATA_reg_RNO[56]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[56]_net_1\, D => 
        \sdr_dataout_reg[8]_net_1\, Y => N_194_mux_i);
    
    \sdr_datain_1[5]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[5]_net_1\, C => \WDATA_reg[53]_net_1\, D
         => \WDATA_reg[37]_net_1\, Y => \sdr_datain_1[5]_net_1\);
    
    \RDATA_reg_RNO[11]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA_0\, D => 
        \sdr_dataout_reg[11]_net_1\, Y => N_181_mux_i);
    
    \sdr_datain_2[6]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[6]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[6]_net_1\);
    
    \WDATA_mux_3_0_0[4]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(4), B => 
        COREAXI_0_AXImslave16_WDATA(36), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[4]_net_1\);
    
    \sdr_datain_0[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[24]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[8]_net_1\);
    
    \WDATA_reg[45]\ : SLE
      port map(D => \WDATA_mux[45]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[45]_net_1\);
    
    un1_sdr_count_0_sqmuxa_0_a2_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \R_VALID\, B => \axi_state[1]_net_1\, Y => 
        N_358);
    
    \WDATA_reg[22]\ : SLE
      port map(D => \WDATA_mux[22]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[22]_net_1\);
    
    \DQM_i_3[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => dqm_sdr, B => \axi_state[0]_net_1\, C => 
        \DQM_mux[1]\, Y => \DQM_i_3[1]_net_1\);
    
    \WDATA_mux_3_0_RNO[13]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[13]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[13]_net_1\, Y => \WDATA_mux_15[13]\);
    
    \RDATA_reg[35]\ : SLE
      port map(D => \sdr_dataout_reg[3]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[35]_net_1\);
    
    OE_xhdl0 : SLE
      port map(D => OE_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => un1_top_sb_0_3_i_i);
    
    \RDATA_reg_RNI1POR[58]\ : CFG4
      generic map(INIT => x"7D41")

      port map(A => \RDATA_reg[58]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        m9_1_1_2, Y => i58_mux);
    
    \asize_reg_RNI8E505[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_6\, C => i22_mux_3_i_1_0, 
        D => i22_mux_3_i_1, Y => i22_mux_3_i);
    
    \asize[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => COREAXI_0_AXImslave16_ARSIZE(0), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWSIZE(0), Y => \asize[0]_net_1\);
    
    \sdr_datain_reg_RNO[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[6]_net_1\, C => \sdr_datain_1[6]_net_1\, Y
         => \sdr_datain[6]\);
    
    \WDATA_reg_RNO[51]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(51), 
        Y => \WDATA_mux[51]\);
    
    axi_nextstate_1_sqmuxa_i_o2_i_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => \N_389\, B => COREAXI_0_AXImslave16_WVALID, C
         => \axi_state[5]_net_1\, Y => \WREADY_SI16\);
    
    \RDATA_reg[51]\ : SLE
      port map(D => N_189_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[51]_net_1\);
    
    \WDATA_mux_8_3[2]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(2), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[2]_net_1\);
    
    \WDATA_reg_RNO[48]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(48), 
        Y => \WDATA_mux[48]\);
    
    \WDATA_mux_3_0_0[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(10), B => 
        COREAXI_0_AXImslave16_WDATA(42), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[10]_net_1\);
    
    \raddr_reg_9_RNO[22]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[22]_net_1\, C => 
        raddr_reg_9_2_axb_22_1, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_21, S => N_771, Y => OPEN, FCO => 
        OPEN);
    
    \axi_state_ns_0[0]\ : CFG4
      generic map(INIT => x"F0F8")

      port map(A => N_23, B => \axi_state_0\, C => 
        \axi_state_ns_0_0[0]_net_1\, D => \N_3297\, Y => 
        \axi_state_ns[0]\);
    
    \WDATA_mux_31[23]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(55), B => 
        COREAXI_0_AXImslave16_WDATA(23), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[23]_net_1\);
    
    \axi_state_ns_0_a2_0[5]\ : CFG4
      generic map(INIT => x"AE00")

      port map(A => \axi_state[5]_net_1\, B => 
        \axi_state[0]_net_1\, C => N_338, D => \N_389\, Y => 
        N_3309);
    
    \WDATA_mux_3_0[4]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[4]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[4]_net_1\, Y => \WDATA_mux[4]\);
    
    \WSTRB_mux_3_0_a3_0_0[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \WSTRB_reg[2]_net_1\, B => 
        \WSTRB_reg[7]_net_1\, Y => 
        \WSTRB_mux_3_0_a3_0_0[3]_net_1\);
    
    \un1_axi_state_4_i_o2_RNIN7N7[0]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_335_i, B => \axi_state[9]_net_1\, Y => 
        raddr_reg_9_sn_N_3_i);
    
    \RDATA_reg[28]\ : SLE
      port map(D => \sdr_dataout_reg[12]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[28]_net_1\);
    
    \WDATA_mux_8_0[4]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(52), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[4]_net_1\);
    
    \WDATA_reg[15]\ : SLE
      port map(D => \WDATA_mux[15]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[15]_net_1\);
    
    \RDATA_reg_RNI5JP32[57]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_3167_i, B => i58_mux_0, Y => 
        COREAXI_0_AXImslave16_RDATA_m_57);
    
    \asize_reg_RNI5B505[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_5\, C => i22_mux_4_i_1_0, 
        D => i22_mux_4_i_1, Y => i22_mux_4_i);
    
    \WDATA_reg[36]\ : SLE
      port map(D => \WDATA_mux[36]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[36]_net_1\);
    
    \sdr_datain_0[6]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[22]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[6]_net_1\);
    
    \sdr_datain_3[9]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[9]_net_1\, C => \WDATA_reg[9]_net_1\, Y => 
        \sdr_datain_3[9]_net_1\);
    
    \WDATA_mux_3_0_RNO[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[6]_net_1\, C => \WDATA_mux_8_1[6]_net_1\, 
        Y => \WDATA_mux_8[6]\);
    
    \sdr_datain_reg_RNO[14]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[14]_net_1\, C => \sdr_datain_1[14]_net_1\, 
        Y => \sdr_datain[14]\);
    
    raddr_reg_9_2_axb_19_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(20), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(20), Y => 
        \raddr_reg_9_2_axb_19_1\);
    
    \WDATA_reg[20]\ : SLE
      port map(D => \WDATA_mux[20]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[20]_net_1\);
    
    \raddr_reg_9[19]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_768, Y => \raddr_reg_9[19]_net_1\);
    
    \WDATA_mux_3_0_0[2]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(2), B => 
        COREAXI_0_AXImslave16_WDATA(34), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[2]_net_1\);
    
    \RDATA_reg_RNO[15]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[15]\, D => 
        \sdr_dataout_reg[15]_net_1\, Y => N_185_mux_i);
    
    \WDATA_reg_RNO[40]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(40), 
        Y => \WDATA_mux[40]\);
    
    \raddr_reg[21]\ : SLE
      port map(D => \raddr_reg_9[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[21]_net_1\);
    
    \raddr_reg_9[14]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_763, Y => \raddr_reg_9[14]_net_1\);
    
    \RDATA_reg_RNIPCDK1[29]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[29]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[13]\, C => N_3141, D => 
        N_3167_i, Y => N_69_mux_i);
    
    \WDATA_mux_3_0_RNO[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[2]_net_1\, C => \WDATA_mux_8_1[2]_net_1\, 
        Y => \WDATA_mux_8[2]\);
    
    \sdr_datain_3[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[2]_net_1\, C => \WDATA_reg[2]_net_1\, Y => 
        \sdr_datain_3[2]_net_1\);
    
    \axi_state_ns_o2[8]\ : CFG4
      generic map(INIT => x"DFFF")

      port map(A => N_71_i, B => un2_sdr_count_NE_0, C => 
        \R_VALID\, D => N_3326_i, Y => N_349);
    
    \WDATA_mux_15_1[12]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[12]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(28), D
         => COREAXI_0_AXImslave16_WDATA(44), Y => 
        \WDATA_mux_15_1[12]_net_1\);
    
    \RDATA_reg_RNI07HJ1[20]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[20]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[4]\, C => N_3141, D => 
        N_3167_i, Y => COREAXI_0_AXImslave16_RDATA_m_20);
    
    \WDATA_mux_3_0_o5[31]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => \N_74\, 
        C => \asize_reg[1]_net_1\, Y => N_3172);
    
    \sdr_datain_reg[6]\ : SLE
      port map(D => \sdr_datain[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(6));
    
    \WDATA_mux_8_0[5]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(53), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[5]_net_1\);
    
    \DQM_i_1[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => dqm_sdr, B => \axi_state[0]_net_1\, C => 
        \DQM_mux[0]\, Y => \DQM_i_1[0]_net_1\);
    
    \WDATA_reg[58]\ : SLE
      port map(D => \WDATA_mux[58]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[58]_net_1\);
    
    \WDATA_reg_RNO[55]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(55), 
        Y => \WDATA_mux[55]\);
    
    \RDATA_reg_RNI6LFQ1[35]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[3]\, B => 
        \RDATA_reg[35]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3169_i);
    
    raddr_reg_9_2_axb_16_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(17), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(17), Y => 
        \raddr_reg_9_2_axb_16_1\);
    
    \axi_state_ns_0_0[7]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => RW_ACK, B => \axi_state[2]_net_1\, C => 
        COREAXI_0_AXImslave16_ARVALID, D => 
        \COREAXI_0_AXImslave16_ARREADY\, Y => 
        \axi_state_ns_0_0[7]_net_1\);
    
    \BA[0]\ : SLE
      port map(D => \BA_i[0]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => BA_c(0));
    
    \RDATA_reg_RNINGEN1[30]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[30]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_0_i_1_0);
    
    \RDATA_reg_RNIIECR1[42]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[10]\, B => 
        \RDATA_reg[42]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_42);
    
    \WDATA_reg[27]\ : SLE
      port map(D => \WDATA_mux[27]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[27]_net_1\);
    
    \sdr_count[2]\ : SLE
      port map(D => N_3278_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_count[2]_net_1\);
    
    \RDATA_reg[18]\ : SLE
      port map(D => N_3071_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[18]_net_1\);
    
    \WDATA_mux_3_0[3]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[3]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[3]_net_1\, Y => \WDATA_mux[3]\);
    
    \RDATA_reg_RNI2UGN1[59]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[59]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_0_i_1);
    
    \WSTRB_mux_8_m1_1[0]\ : CFG4
      generic map(INIT => x"10DC")

      port map(A => \WSTRB_reg[5]_net_1\, B => 
        \WSTRB_reg[4]_net_1\, C => \WSTRB_reg[6]_net_1\, D => 
        \WSTRB_reg[3]_net_1\, Y => \WSTRB_mux_8_m1_1[0]_net_1\);
    
    \axi_state_ns_i_a2[4]\ : CFG4
      generic map(INIT => x"0301")

      port map(A => \axi_state[0]_net_1\, B => 
        \COREAXI_0_AXImslave16_AWREADY\, C => 
        \axi_state[5]_net_1\, D => N_338, Y => N_368);
    
    \WDATA_mux_3[21]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(21), C => 
        \WDATA_mux_31[21]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[21]\);
    
    \raddr_reg_RNIOKL3I[12]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[12]_net_1\, C => 
        \raddr_reg_9_2_axb_12_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_11, S => N_761, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_12);
    
    \sdr_dataout_reg[1]\ : SLE
      port map(D => DQ_in(1), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[1]_net_1\);
    
    \axi_state[0]\ : SLE
      port map(D => \axi_state_ns[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[0]_net_1\);
    
    \raddr_reg[11]\ : SLE
      port map(D => \raddr_reg_9[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[11]_net_1\);
    
    \DQM[0]\ : SLE
      port map(D => \DQM_i_1[0]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        DQM_c(0));
    
    \sdr_datain_0[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[18]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[2]_net_1\);
    
    \WDATA_mux_31[22]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(54), B => 
        COREAXI_0_AXImslave16_WDATA(22), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[22]_net_1\);
    
    \WDATA_reg[24]\ : SLE
      port map(D => \WDATA_mux[24]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[24]_net_1\);
    
    \RDATA_reg_RNINETB1[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[2]\, Y => N_39);
    
    \WDATA_mux_8_0[6]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(54), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[6]_net_1\);
    
    \un7_1.SUM_i_o2[3]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \COREAXI_0_AXImslave16_ARREADY\, B => 
        \axi_state[9]_net_1\, C => 
        \COREAXI_0_AXImslave16_AWREADY\, D => 
        \COREAXI_0_AXImslave16_BVALID\, Y => N_3293);
    
    \raddr_reg_9_2_1_1[1]\ : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(2), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(2), Y => 
        \raddr_reg_9_2_1_1[1]_net_1\);
    
    \DQM_mux_ns_1_1[0]\ : CFG3
      generic map(INIT => x"1D")

      port map(A => \WSTRB_reg[4]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \WSTRB_reg[6]_net_1\, Y => 
        \DQM_mux_ns_1_1[0]_net_1\);
    
    \RDATA_reg_RNI29HJ1[21]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[21]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[5]\, C => N_3141, D => 
        N_3167_i, Y => COREAXI_0_AXImslave16_RDATA_m_21);
    
    \WDATA_mux_3_0_0[12]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(12), B => 
        COREAXI_0_AXImslave16_WDATA(44), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[12]_net_1\);
    
    \RDATA_reg[41]\ : SLE
      port map(D => \sdr_dataout_reg[9]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[41]_net_1\);
    
    \WDATA_mux_8_3[5]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(5), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[5]_net_1\);
    
    \sdr_datain_reg[11]\ : SLE
      port map(D => \sdr_datain[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(11));
    
    \sdr_datain_0[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[16]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[0]_net_1\);
    
    \WDATA_reg[39]\ : SLE
      port map(D => \WDATA_mux[39]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[39]_net_1\);
    
    \RDATA_reg_RNO[7]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[7]\, D => 
        \sdr_dataout_reg[7]_net_1\, Y => N_177_mux_i);
    
    raddr_reg_9_2_axb_7_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(8), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(8), Y => 
        \raddr_reg_9_2_axb_7_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \WDATA_reg_RNO[62]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(62), 
        Y => \WDATA_mux[62]\);
    
    \raddr_reg[17]\ : SLE
      port map(D => \raddr_reg_9[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[17]_net_1\);
    
    \RDATA_reg_RNIETFQ1[39]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[7]\, B => 
        \RDATA_reg[39]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3096_i);
    
    \WDATA_reg_RNO[46]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(46), 
        Y => \WDATA_mux[46]\);
    
    \SA[2]\ : SLE
      port map(D => \SA_i[2]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(2));
    
    raddr_reg_9_2_axb_4_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(5), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(5), Y => 
        \raddr_reg_9_2_axb_4_1\);
    
    \raddr_reg_9[1]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_750, Y => \raddr_reg_9[1]_net_1\);
    
    \WDATA_reg[6]\ : SLE
      port map(D => \WDATA_mux[6]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[6]_net_1\);
    
    \RDATA_reg[5]\ : SLE
      port map(D => N_175_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[5]\);
    
    \axi_count[3]\ : SLE
      port map(D => N_3271_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_count[3]_net_1\);
    
    \WDATA_mux_3_0[16]\ : CFG4
      generic map(INIT => x"CECC")

      port map(A => N_3157, B => \WDATA_mux_3_0_0[16]_net_1\, C
         => COREAXI_0_AXImslave16_WSTRB(2), D => 
        \WDATA_mux_8_m0[0]\, Y => \WDATA_mux[16]\);
    
    \raddr_reg_RNIGVTDA[6]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[6]_net_1\, C => 
        \raddr_reg_9_2_axb_6_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_5, S => N_755, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_6);
    
    \RDATA_reg_RNO[14]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA_3\, D => 
        \sdr_dataout_reg[14]_net_1\, Y => N_184_mux_i);
    
    \WDATA_mux_3_0_RNO[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[0]_net_1\, C => \WDATA_mux_8_1[0]_net_1\, 
        Y => \WDATA_mux_8[0]\);
    
    \WDATA_mux_3_0_m4[15]\ : CFG3
      generic map(INIT => x"AD")

      port map(A => \asize_reg[1]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => \asize_reg[0]_net_1\, 
        Y => N_3210);
    
    raddr_reg_9_2_axb_14_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(15), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(15), Y => 
        \raddr_reg_9_2_axb_14_1\);
    
    \sdr_datain_1[2]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[2]_net_1\, C => \WDATA_reg[50]_net_1\, D
         => \WDATA_reg[34]_net_1\, Y => \sdr_datain_1[2]_net_1\);
    
    \sdr_count_RNIQ0CH1[3]\ : CFG4
      generic map(INIT => x"5556")

      port map(A => \sdr_count[3]_net_1\, B => 
        \B_SIZE_reg[2]_net_1\, C => \B_SIZE_reg[1]_net_1\, D => 
        \B_SIZE_reg[0]_net_1\, Y => N_71_i);
    
    \axi_count_7_i_o2_1[0]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \axi_count[0]_net_1\, B => 
        \COREAXI_0_AXImslave16_AWREADY\, C => 
        \COREAXI_0_AXImslave16_ARREADY\, Y => N_72);
    
    \raddr_reg[20]\ : SLE
      port map(D => \raddr_reg_9[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[20]_net_1\);
    
    \RDATA_reg_RNIF9L42[58]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_3167_i, B => i58_mux, Y => 
        COREAXI_0_AXImslave16_RDATA_m_58);
    
    \RDATA_reg_RNI4BHJ1[22]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[22]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[6]\, C => N_3141, D => 
        N_3167_i, Y => N_80_mux_i);
    
    \WDATA_mux_8_0[1]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(49), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[1]_net_1\);
    
    \WDATA_mux_3_0_a5_0[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => COREAXI_0_AXImslave16_WSTRB(1), B => 
        COREAXI_0_AXImslave16_WDATA(14), C => 
        \asize_reg[1]_net_1\, Y => N_3200);
    
    \WDATA_mux_3_0_0[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(6), B => 
        COREAXI_0_AXImslave16_WDATA(38), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[6]_net_1\);
    
    \WDATA_mux_3_0[15]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[15]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[15]_net_1\, Y => \WDATA_mux[15]\);
    
    \raddr_reg[14]\ : SLE
      port map(D => \raddr_reg_9[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[14]_net_1\);
    
    \WDATA_reg_RNO[32]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(32), 
        Y => \WDATA_mux[32]\);
    
    \axi_state_ns_o2[9]\ : CFG4
      generic map(INIT => x"DFFF")

      port map(A => N_71_i, B => un2_sdr_count_NE_0, C => W_VALID, 
        D => N_3326_i, Y => N_338);
    
    \un1_B_SIZE_reg_0_a2[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \B_SIZE_reg[1]_net_1\, B => N_335_i, C => 
        N_343_i, Y => \un1_B_SIZE_reg_0_a2[1]_net_1\);
    
    \WDATA_mux_8_1[1]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[1]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(33), D
         => COREAXI_0_AXImslave16_WDATA(17), Y => 
        \WDATA_mux_8_1[1]_net_1\);
    
    \sdr_datain_3[1]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[1]_net_1\, C => \WDATA_reg[1]_net_1\, Y => 
        \sdr_datain_3[1]_net_1\);
    
    \WDATA_reg_RNO[54]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(54), 
        Y => \WDATA_mux[54]\);
    
    \sdr_count_RNO[2]\ : CFG4
      generic map(INIT => x"0041")

      port map(A => N_3281, B => N_3288, C => 
        \sdr_count[2]_net_1\, D => N_3293, Y => N_3278_i);
    
    \RDATA_reg_RNO[8]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[8]\, D => 
        \sdr_dataout_reg[8]_net_1\, Y => N_178_mux_i);
    
    raddr_reg_9_2_axb_11_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(12), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(12), Y => 
        \raddr_reg_9_2_axb_11_1\);
    
    \raddr_reg[22]\ : SLE
      port map(D => \raddr_reg_9[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[22]_net_1\);
    
    \WDATA_mux_15_0[13]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(61), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[13]_net_1\);
    
    \RDATA_reg[23]\ : SLE
      port map(D => \sdr_dataout_reg[7]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[23]_net_1\);
    
    \raddr_reg_9[0]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => \un1_B_SIZE_reg_0_a2_RNISOQQ1_Y[2]\, Y => 
        \raddr_reg_9[0]_net_1\);
    
    \SA[0]\ : SLE
      port map(D => \SA_i[0]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(0));
    
    \WDATA_reg[41]\ : SLE
      port map(D => \WDATA_mux[41]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[41]_net_1\);
    
    \WDATA_mux_31[20]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(52), B => 
        COREAXI_0_AXImslave16_WDATA(20), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[20]_net_1\);
    
    \RDATA_reg_RNO[53]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[53]_net_1\, D => 
        \sdr_dataout_reg[5]_net_1\, Y => N_191_mux_i);
    
    \RDATA_reg_RNIBFPC1[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[15]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_15\);
    
    \WDATA_reg[35]\ : SLE
      port map(D => \WDATA_mux[35]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[35]_net_1\);
    
    \BA[1]\ : SLE
      port map(D => \BA_i[1]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => BA_c(1));
    
    \RDATA_reg[31]\ : SLE
      port map(D => N_3074_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[31]_net_1\);
    
    \RDATA_reg_RNI0FFQ1[32]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[0]\, B => 
        \RDATA_reg[32]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3066_i);
    
    \raddr_reg[10]\ : SLE
      port map(D => \raddr_reg_9[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[10]_net_1\);
    
    \RDATA_reg_RNILCTB1[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[0]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_0\);
    
    \RDATA_reg_RNIQHTB1[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[5]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_5\);
    
    \RDATA_reg_RNINADK1[28]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[28]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[12]\, C => N_3141, D => 
        N_3167_i, Y => N_75_mux_i);
    
    \WSTRB_mux_3_0_m3[0]\ : CFG4
      generic map(INIT => x"AAAC")

      port map(A => \WSTRB_reg[0]_net_1\, B => 
        \WSTRB_mux_8_m1[0]_net_1\, C => N_3141, D => N_26, Y => 
        N_3145);
    
    \sdr_datain_3[8]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[8]_net_1\, C => \WDATA_reg[8]_net_1\, Y => 
        \sdr_datain_3[8]_net_1\);
    
    \RDATA_reg_RNISOHN1[62]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[62]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_0_i_1);
    
    \WDATA_reg[26]\ : SLE
      port map(D => \WDATA_mux[26]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[26]_net_1\);
    
    \axi_state[2]\ : SLE
      port map(D => \axi_state_ns[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[2]_net_1\);
    
    \CS_N[0]\ : SLE
      port map(D => \CS_N_i[0]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => CS_N_c_0);
    
    \RDATA_reg[62]\ : SLE
      port map(D => N_200_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[62]_net_1\);
    
    \asize_reg_RNIOC315[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_15\, C => i17_mux_i_1_0, D
         => i17_mux_i_1, Y => i17_mux_i);
    
    \axi_count[1]\ : SLE
      port map(D => N_3273_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_count[1]_net_1\);
    
    \raddr_reg[7]\ : SLE
      port map(D => \raddr_reg_9[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[7]_net_1\);
    
    \raddr_reg[12]\ : SLE
      port map(D => \raddr_reg_9[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[12]_net_1\);
    
    \WDATA_reg[53]\ : SLE
      port map(D => \WDATA_mux[53]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[53]_net_1\);
    
    \WDATA_mux_8_3[6]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(6), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[6]_net_1\);
    
    \WDATA_reg[11]\ : SLE
      port map(D => \WDATA_mux[11]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[11]_net_1\);
    
    \RDATA_reg[58]\ : SLE
      port map(D => N_196_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[58]_net_1\);
    
    \WDATA_mux_3[18]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(18), C => 
        \WDATA_mux_31[18]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[18]\);
    
    \WDATA_mux_8_0[3]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(51), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[3]_net_1\);
    
    \WDATA_mux_3_0[12]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[12]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[12]_net_1\, Y => \WDATA_mux[12]\);
    
    \WSTRB_mux_8_m1_1[1]\ : CFG4
      generic map(INIT => x"10BA")

      port map(A => \WSTRB_reg[5]_net_1\, B => 
        \WSTRB_reg[4]_net_1\, C => \WSTRB_reg[7]_net_1\, D => 
        \WSTRB_reg[2]_net_1\, Y => \WSTRB_mux_8_m1_1[1]_net_1\);
    
    \raddr_reg[8]\ : SLE
      port map(D => \raddr_reg_9[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[8]_net_1\);
    
    \WDATA_reg[8]\ : SLE
      port map(D => \WDATA_mux[8]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[8]_net_1\);
    
    \RDATA_reg_RNIP5O32[50]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_3167_i, B => i58_mux_1, Y => 
        COREAXI_0_AXImslave16_RDATA_m_50);
    
    \WDATA_reg[63]\ : SLE
      port map(D => \WDATA_mux[63]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[63]_net_1\);
    
    \axi_state_ns_0_0[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_BVALID, B => 
        N_3313, C => \COREAXI_0_AXImslave16_BVALID\, Y => 
        \axi_state_ns_0_0[0]_net_1\);
    
    \RDATA_reg_RNO[59]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[59]_net_1\, D => 
        \sdr_dataout_reg[11]_net_1\, Y => N_197_mux_i);
    
    \RDATA_reg_RNIRITB1[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[6]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_6\);
    
    \RDATA_reg[13]\ : SLE
      port map(D => N_183_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[13]\);
    
    \raddr_reg_RNIRNRN6[3]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[3]_net_1\, C => 
        \raddr_reg_9_2_axb_3_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_2, S => N_752, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_3);
    
    \raddr_reg_RNI6FI69[5]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[5]_net_1\, C => 
        \raddr_reg_9_2_axb_5_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_4, S => N_754, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_5);
    
    \WDATA_reg[3]\ : SLE
      port map(D => \WDATA_mux[3]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[3]_net_1\);
    
    \sdr_datain_reg_RNO[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[13]_net_1\, C => \sdr_datain_1[13]_net_1\, 
        Y => \sdr_datain[13]\);
    
    \SA[10]\ : SLE
      port map(D => \SA_i[10]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(10));
    
    \raddr_reg[5]\ : SLE
      port map(D => \raddr_reg_9[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[5]_net_1\);
    
    \sdr_datain_reg[8]\ : SLE
      port map(D => \sdr_datain[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(8));
    
    \RDATA_reg_RNI0H7C[18]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \COREAXI_0_AXImslave16_RDATA[2]\, B => 
        \asize_reg[0]_net_1\, C => \RDATA_reg[18]_net_1\, Y => 
        m23_1_2);
    
    un5_axi_rvalid_i_0_o2 : CFG2
      generic map(INIT => x"7")

      port map(A => COREAXI_0_AXImslave16_ARVALID, B => 
        COREAXI_0_AXImslave16_ARBURST_0, Y => un5_axi_rvalid_i_0);
    
    \RDATA_reg[7]\ : SLE
      port map(D => N_177_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[7]\);
    
    \sdr_datain_0[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[25]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[9]_net_1\);
    
    \axi_state[7]\ : SLE
      port map(D => \axi_state_ns[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_AWREADY\);
    
    \raddr_reg_9_2_1_1[2]\ : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(3), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(3), Y => 
        \raddr_reg_9_2_1_1[2]_net_1\);
    
    \sdr_datain_2[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[15]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[15]_net_1\);
    
    \sdr_datain_reg_RNO[15]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[15]_net_1\, C => \sdr_datain_1[15]_net_1\, 
        Y => \sdr_datain[15]\);
    
    \WDATA_mux_15_0[14]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(62), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[14]_net_1\);
    
    \WSTRB_reg[4]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(4), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[4]_net_1\);
    
    \raddr_reg_RNIOTA71[0]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => \raddr_reg[0]_net_1\, B => 
        \raddr_reg_9_2_1_1[0]_net_1\, C => raddr_reg_9_sn_N_3_i, 
        Y => \raddr_reg_RNIOTA71[0]_net_1\);
    
    \raddr_reg_9[18]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_767, Y => \raddr_reg_9[18]_net_1\);
    
    \RDATA_reg[60]\ : SLE
      port map(D => N_198_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[60]_net_1\);
    
    \WDATA_reg[1]\ : SLE
      port map(D => \WDATA_mux[1]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[1]_net_1\);
    
    \RDATA_reg_RNI0RFN1[48]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[48]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_2_i_1);
    
    \raddr_reg[18]\ : SLE
      port map(D => \raddr_reg_9[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[18]_net_1\);
    
    \sdr_datain_reg_RNO[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[2]_net_1\, C => \sdr_datain_1[2]_net_1\, Y
         => \sdr_datain[2]\);
    
    \WDATA_reg_RNO[38]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(38), 
        Y => \WDATA_mux[38]\);
    
    \WDATA_mux_3_0[14]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => \asize_reg[0]_net_1\, B => 
        \asize_reg[1]_net_1\, C => \WDATA_mux_3_0_1[14]_net_1\, D
         => \WDATA_mux_15[14]\, Y => \WDATA_mux[14]\);
    
    \sdr_datain_reg[5]\ : SLE
      port map(D => \sdr_datain[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(5));
    
    \RDATA_reg_RNO[31]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[31]_net_1\, D => 
        \sdr_dataout_reg[15]_net_1\, Y => N_3074_i);
    
    \RDATA_reg_RNI5N8C[25]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \COREAXI_0_AXImslave16_RDATA[9]\, B => 
        \asize_reg[0]_net_1\, C => \RDATA_reg[25]_net_1\, Y => 
        m16_1_1_2);
    
    \RDATA_reg_RNIAHHJ1[25]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[25]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[9]\, C => N_3141, D => 
        N_3167_i, Y => N_78_mux_i);
    
    raddr_reg_9_2_axb_12_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(13), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(13), Y => 
        \raddr_reg_9_2_axb_12_1\);
    
    \WDATA_reg_RNO[60]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(60), 
        Y => \WDATA_mux[60]\);
    
    \WDATA_reg[29]\ : SLE
      port map(D => \WDATA_mux[29]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[29]_net_1\);
    
    \sdr_datain_reg[3]\ : SLE
      port map(D => \sdr_datain[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(3));
    
    \un1_B_SIZE_reg_0_a2_RNIQJLL3[1]\ : ARI1
      generic map(INIT => x"5758A")

      port map(A => \raddr_reg_RNIR0B71[1]_net_1\, B => 
        \un1_B_SIZE_reg_0_a2[1]_net_1\, C => N_335_i, D => 
        \axi_state[9]_net_1\, FCI => raddr_reg_9_2_cry_0, S => 
        N_750, Y => OPEN, FCO => raddr_reg_9_2_cry_1);
    
    \WSTRB_mux_8_m1[1]\ : CFG4
      generic map(INIT => x"FAF8")

      port map(A => \WSTRB_mux_8_m1_1[1]_net_1\, B => 
        \un7_wstrb_reg_i_a3\, C => \WSTRB_reg[3]_net_1\, D => 
        \WSTRB_reg[5]_net_1\, Y => \WSTRB_mux_8_m1[1]_net_1\);
    
    \sdr_datain_2[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[12]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[12]_net_1\);
    
    \raddr_reg_RNIQ12UO[17]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[17]_net_1\, C => 
        \raddr_reg_9_2_axb_17_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_16, S => N_766, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_17);
    
    \WDATA_mux_8_1[2]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[2]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(34), D
         => COREAXI_0_AXImslave16_WDATA(18), Y => 
        \WDATA_mux_8_1[2]_net_1\);
    
    \sdr_datain_2[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[2]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[2]_net_1\);
    
    \SA[1]\ : SLE
      port map(D => \SA_i[1]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(1));
    
    \WDATA_mux_15_3[13]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(13), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[13]_net_1\);
    
    \asize_reg_RNIL9315[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_14\, C => i17_mux_0_i_1_0, 
        D => i17_mux_0_i_1, Y => i17_mux_0_i);
    
    \sdr_dataout_reg[5]\ : SLE
      port map(D => DQ_in(5), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[5]_net_1\);
    
    \raddr_reg_RNIR0B71[1]\ : CFG4
      generic map(INIT => x"B1F0")

      port map(A => N_335_i, B => \raddr_reg_9_2_1_1[1]_net_1\, C
         => \raddr_reg[1]_net_1\, D => \axi_state[9]_net_1\, Y
         => \raddr_reg_RNIR0B71[1]_net_1\);
    
    \RDATA_reg_RNO[2]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[2]\, D => 
        \sdr_dataout_reg[2]_net_1\, Y => N_172_mux_i);
    
    \WDATA_mux_8_3[4]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(4), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[4]_net_1\);
    
    \WSTRB_mux_3_0_a3[1]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \WSTRB_reg[0]_net_1\, B => 
        \WSTRB_reg[5]_net_1\, C => \un7_wstrb_reg_i_a3\, D => 
        N_3157, Y => N_3153);
    
    \sdr_datain_1[8]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[8]_net_1\, C => \WDATA_reg[56]_net_1\, D
         => \WDATA_reg[40]_net_1\, Y => \sdr_datain_1[8]_net_1\);
    
    \RDATA_reg_RNIULTB1[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[9]\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_9);
    
    \sdr_dataout_reg[13]\ : SLE
      port map(D => DQ_in(13), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[13]_net_1\);
    
    \RDATA_reg[9]\ : SLE
      port map(D => N_179_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[9]\);
    
    \sdr_count[1]\ : SLE
      port map(D => N_3279_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_count[1]_net_1\);
    
    \un1_B_SIZE_reg_0_a2[0]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \B_SIZE_reg[2]_net_1\, B => N_335_i, C => 
        N_343_i, Y => \un1_B_SIZE_reg_0_a2[0]_net_1\);
    
    \WDATA_mux_15_0[15]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(63), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[15]_net_1\);
    
    \RDATA_reg_RNIRMGN1[52]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[52]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_5_i_1);
    
    \axi_state[6]\ : SLE
      port map(D => \axi_state_ns[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state_0\);
    
    \raddr_reg[9]\ : SLE
      port map(D => \raddr_reg_9[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[9]_net_1\);
    
    \raddr_reg_RNIPUACF[10]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[10]_net_1\, C => 
        \raddr_reg_9_2_axb_10_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_9, S => N_759, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_10);
    
    \RDATA_reg_RNIPHDN1[23]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[23]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_2_i_1_0);
    
    \raddr_reg_RNIT0O9Q[18]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[18]_net_1\, C => 
        \raddr_reg_9_2_axb_18_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_17, S => N_767, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_18);
    
    \WDATA_reg_RNO[43]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(43), 
        Y => \WDATA_mux[43]\);
    
    \axi_state_RNI5FHE[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => COREAXI_0_AXImslave16_WVALID, B => 
        \axi_state[5]_net_1\, C => \axi_state[3]_net_1\, Y => 
        N_355_i);
    
    \RDATA_reg[48]\ : SLE
      port map(D => N_186_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[48]_net_1\);
    
    \WDATA_mux_15_0[9]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(57), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[9]_net_1\);
    
    \RDATA_reg_RNIJ6DK1[26]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[26]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[10]\, C => N_3141, D => 
        N_3167_i, Y => N_77_mux_i);
    
    \RDATA_reg_RNI8CPC1[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[12]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_12\);
    
    \WDATA_mux_3_0_a4_0[31]\ : CFG3
      generic map(INIT => x"40")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => N_3157, 
        C => COREAXI_0_AXImslave16_WSTRB(7), Y => N_3207);
    
    \RDATA_reg_RNITLDN1[27]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[27]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_0_i_1_0);
    
    CoreSDR_0 : CORESDR
      port map(RADDR(30) => GND_net_1, RADDR(29) => GND_net_1, 
        RADDR(28) => GND_net_1, RADDR(27) => GND_net_1, RADDR(26)
         => GND_net_1, RADDR(25) => GND_net_1, RADDR(24) => 
        GND_net_1, RADDR(23) => GND_net_1, RADDR(22) => 
        \raddr_reg[22]_net_1\, RADDR(21) => \raddr_reg[21]_net_1\, 
        RADDR(20) => \raddr_reg[20]_net_1\, RADDR(19) => 
        \raddr_reg[19]_net_1\, RADDR(18) => \raddr_reg[18]_net_1\, 
        RADDR(17) => \raddr_reg[17]_net_1\, RADDR(16) => 
        \raddr_reg[16]_net_1\, RADDR(15) => \raddr_reg[15]_net_1\, 
        RADDR(14) => \raddr_reg[14]_net_1\, RADDR(13) => 
        \raddr_reg[13]_net_1\, RADDR(12) => \raddr_reg[12]_net_1\, 
        RADDR(11) => \raddr_reg[11]_net_1\, RADDR(10) => 
        \raddr_reg[10]_net_1\, RADDR(9) => \raddr_reg[9]_net_1\, 
        RADDR(8) => \raddr_reg[8]_net_1\, RADDR(7) => 
        \raddr_reg[7]_net_1\, RADDR(6) => \raddr_reg[6]_net_1\, 
        RADDR(5) => \raddr_reg[5]_net_1\, RADDR(4) => 
        \raddr_reg[4]_net_1\, RADDR(3) => \raddr_reg[3]_net_1\, 
        RADDR(2) => \raddr_reg[2]_net_1\, RADDR(1) => 
        \raddr_reg[1]_net_1\, RADDR(0) => \raddr_reg[0]_net_1\, 
        B_SIZE(3) => GND_net_1, B_SIZE(2) => 
        \B_SIZE_reg[2]_net_1\, B_SIZE(1) => \B_SIZE_reg[1]_net_1\, 
        B_SIZE(0) => \B_SIZE_reg[0]_net_1\, RAS(3) => GND_net_1, 
        RAS(2) => GND_net_1, RAS(1) => VCC_net_1, RAS(0) => 
        GND_net_1, RCD(2) => GND_net_1, RCD(1) => VCC_net_1, 
        RCD(0) => GND_net_1, RRD(1) => VCC_net_1, RRD(0) => 
        GND_net_1, RP(2) => GND_net_1, RP(1) => VCC_net_1, RP(0)
         => VCC_net_1, RC(3) => VCC_net_1, RC(2) => GND_net_1, 
        RC(1) => GND_net_1, RC(0) => GND_net_1, RFC(3) => 
        VCC_net_1, RFC(2) => GND_net_1, RFC(1) => GND_net_1, 
        RFC(0) => VCC_net_1, WR(1) => VCC_net_1, WR(0) => 
        GND_net_1, MRD(2) => GND_net_1, MRD(1) => VCC_net_1, 
        MRD(0) => GND_net_1, CL(2) => GND_net_1, CL(1) => 
        VCC_net_1, CL(0) => GND_net_1, BL(1) => VCC_net_1, BL(0)
         => VCC_net_1, DELAY(15) => GND_net_1, DELAY(14) => 
        GND_net_1, DELAY(13) => GND_net_1, DELAY(12) => VCC_net_1, 
        DELAY(11) => VCC_net_1, DELAY(10) => GND_net_1, DELAY(9)
         => VCC_net_1, DELAY(8) => GND_net_1, DELAY(7) => 
        VCC_net_1, DELAY(6) => GND_net_1, DELAY(5) => GND_net_1, 
        DELAY(4) => VCC_net_1, DELAY(3) => GND_net_1, DELAY(2)
         => GND_net_1, DELAY(1) => GND_net_1, DELAY(0) => 
        GND_net_1, REF(15) => GND_net_1, REF(14) => GND_net_1, 
        REF(13) => GND_net_1, REF(12) => VCC_net_1, REF(11) => 
        GND_net_1, REF(10) => GND_net_1, REF(9) => GND_net_1, 
        REF(8) => GND_net_1, REF(7) => GND_net_1, REF(6) => 
        GND_net_1, REF(5) => GND_net_1, REF(4) => GND_net_1, 
        REF(3) => GND_net_1, REF(2) => GND_net_1, REF(1) => 
        GND_net_1, REF(0) => GND_net_1, COLBITS(2) => GND_net_1, 
        COLBITS(1) => VCC_net_1, COLBITS(0) => VCC_net_1, 
        ROWBITS(1) => GND_net_1, ROWBITS(0) => VCC_net_1, SA(13)
         => nc2, SA(12) => nc1, SA(11) => \SA_i[11]\, SA(10) => 
        \SA_i[10]\, SA(9) => \SA_i[9]\, SA(8) => \SA_i[8]\, SA(7)
         => \SA_i[7]\, SA(6) => \SA_i[6]\, SA(5) => \SA_i[5]\, 
        SA(4) => \SA_i[4]\, SA(3) => \SA_i[3]\, SA(2) => 
        \SA_i[2]\, SA(1) => \SA_i[1]\, SA(0) => \SA_i[0]\, BA(1)
         => \BA_i[1]\, BA(0) => \BA_i[0]\, CS_N(0) => \CS_N_i[0]\, 
        CLK => SDRCLK_c, RESET_N => MSS_READY, R_REQ => 
        \un3_r_req_0_0\, W_REQ => N_355_i, AUTO_PCH => GND_net_1, 
        SD_INIT => GND_net_1, REGDIMM => GND_net_1, RW_ACK => 
        RW_ACK, R_VALID => R_VALID_i, D_REQ => OPEN, W_VALID => 
        W_VALID, OE => OE_i, DQM => dqm_sdr, CKE => CKE_i, RAS_N
         => RAS_N_i, CAS_N => CAS_N_i, WE_N => WE_N_i);
    
    \RDATA_reg_RNO[17]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[17]_net_1\, D => 
        \sdr_dataout_reg[1]_net_1\, Y => N_3070_i);
    
    \un7_1.N_3273_i\ : CFG3
      generic map(INIT => x"09")

      port map(A => N_3289, B => \axi_count[1]_net_1\, C => 
        N_3293, Y => N_3273_i);
    
    \RDATA_reg_RNO[48]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[48]_net_1\, D => 
        \sdr_dataout_reg[0]_net_1\, Y => N_186_mux_i);
    
    \WDATA_mux_8_3[7]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(7), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[7]_net_1\);
    
    \WDATA_mux_31[19]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(51), B => 
        COREAXI_0_AXImslave16_WDATA(19), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[19]_net_1\);
    
    \WDATA_reg[25]\ : SLE
      port map(D => \WDATA_mux[25]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[25]_net_1\);
    
    \DQM_mux_ns_1[0]\ : CFG4
      generic map(INIT => x"5702")

      port map(A => \sdr_count[1]_net_1\, B => 
        \DQM_mux_ns_1_1[0]_net_1\, C => \N_74\, D => 
        \WSTRB_mux[2]\, Y => \DQM_mux_ns_1[0]_net_1\);
    
    \sdr_count_RNIPVBH1[2]\ : CFG4
      generic map(INIT => x"9996")

      port map(A => \sdr_count[2]_net_1\, B => 
        \B_SIZE_reg[2]_net_1\, C => \B_SIZE_reg[1]_net_1\, D => 
        \B_SIZE_reg[0]_net_1\, Y => N_3326_i);
    
    \WSTRB_reg[2]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(2), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[2]_net_1\);
    
    \sdr_datain_reg_RNO[11]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[11]_net_1\, C => \sdr_datain_1[11]_net_1\, 
        Y => \sdr_datain[11]\);
    
    \sdr_count_9_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_3281, B => N_3293, Y => N_3299);
    
    \WDATA_reg_RNO[57]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(57), 
        Y => \WDATA_mux[57]\);
    
    \sdr_datain_3[15]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[15]_net_1\, C => \WDATA_reg[15]_net_1\, Y
         => \sdr_datain_3[15]_net_1\);
    
    \RDATA_reg_RNO[51]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[51]_net_1\, D => 
        \sdr_dataout_reg[3]_net_1\, Y => N_189_mux_i);
    
    \asize_reg_RNIF2JA[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \asize_reg[1]_net_1\, B => 
        \asize_reg[0]_net_1\, Y => \N_74\);
    
    \WDATA_mux_15_3[9]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(9), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[9]_net_1\);
    
    \sdr_dataout_reg[7]\ : SLE
      port map(D => DQ_in(7), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[7]_net_1\);
    
    \sdr_datain_2[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[9]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[9]_net_1\);
    
    \RDATA_reg_RNIQIDN1[24]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[24]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_1_i_1_0);
    
    \WDATA_mux_3_0_RNO[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[3]_net_1\, C => \WDATA_mux_8_1[3]_net_1\, 
        Y => \WDATA_mux_8[3]\);
    
    \RDATA_reg[1]\ : SLE
      port map(D => N_171_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[1]\);
    
    \RDATA_reg_RNO[62]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[62]_net_1\, D => 
        \sdr_dataout_reg[14]_net_1\, Y => N_200_mux_i);
    
    \RDATA_reg_RNI7DGJ1[19]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[19]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[3]\, C => N_3141, D => 
        N_3167_i, Y => COREAXI_0_AXImslave16_RDATA_m_19);
    
    \raddr_reg_9[17]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_766, Y => \raddr_reg_9[17]_net_1\);
    
    \WDATA_mux_8_1[3]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[3]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(35), D
         => COREAXI_0_AXImslave16_WDATA(19), Y => 
        \WDATA_mux_8_1[3]_net_1\);
    
    \RDATA_reg[53]\ : SLE
      port map(D => N_191_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[53]_net_1\);
    
    \WDATA_mux_3_0_1[14]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => COREAXI_0_AXImslave16_WDATA(14), B => N_3200, 
        C => \N_74\, D => N_3202, Y => 
        \WDATA_mux_3_0_1[14]_net_1\);
    
    \WDATA_mux_3_0[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(59), B => 
        COREAXI_0_AXImslave16_WDATA(27), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[27]\);
    
    \RDATA_reg[8]\ : SLE
      port map(D => N_178_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[8]\);
    
    \WDATA_reg_RNO[49]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(49), 
        Y => \WDATA_mux[49]\);
    
    \WDATA_reg[31]\ : SLE
      port map(D => \WDATA_mux[31]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[31]_net_1\);
    
    \raddr_reg_9[7]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_756, Y => \raddr_reg_9[7]_net_1\);
    
    \WDATA_mux_15_3[14]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(14), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[14]_net_1\);
    
    \sdr_datain_reg_RNO[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[5]_net_1\, C => \sdr_datain_1[5]_net_1\, Y
         => \sdr_datain[5]\);
    
    \WSTRB_mux_3_0[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \WSTRB_reg[2]_net_1\, B => 
        \WSTRB_mux_3_0_a3_0_0[2]_net_1\, C => N_3149_2, D => 
        N_3141, Y => \WSTRB_mux[2]\);
    
    \sdr_dataout_reg[12]\ : SLE
      port map(D => DQ_in(12), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[12]_net_1\);
    
    \sdr_datain_1[3]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[3]_net_1\, C => \WDATA_reg[51]_net_1\, D
         => \WDATA_reg[35]_net_1\, Y => \sdr_datain_1[3]_net_1\);
    
    \RDATA_reg_RNIRNHN1[61]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[61]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_1_i_1);
    
    \sdr_datain_3[12]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[12]_net_1\, C => \WDATA_reg[12]_net_1\, Y
         => \sdr_datain_3[12]_net_1\);
    
    \WDATA_reg_RNO[36]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(36), 
        Y => \WDATA_mux[36]\);
    
    \WDATA_mux_3_0_RNO[8]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[8]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[8]_net_1\, Y => \WDATA_mux_15[8]\);
    
    \raddr_reg_9[22]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_771, Y => \raddr_reg_9[22]_net_1\);
    
    \WDATA_reg[48]\ : SLE
      port map(D => \WDATA_mux[48]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[48]_net_1\);
    
    \WDATA_mux_3_0[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[1]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[1]_net_1\, Y => \WDATA_mux[1]\);
    
    \RDATA_reg_RNIAEPC1[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA_3\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_14\);
    
    \RDATA_reg_RNIPGTB1[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[4]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_4\);
    
    \RDATA_reg[38]\ : SLE
      port map(D => \sdr_dataout_reg[6]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[38]_net_1\);
    
    \raddr_reg_9[2]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_751, Y => \raddr_reg_9[2]_net_1\);
    
    \RDATA_reg[22]\ : SLE
      port map(D => \sdr_dataout_reg[6]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[22]_net_1\);
    
    \SA[11]\ : SLE
      port map(D => \SA_i[11]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(11));
    
    \RDATA_reg_RNI7BPC1[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA_0\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_11\);
    
    \RDATA_reg_RNIUE7C[17]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \COREAXI_0_AXImslave16_RDATA[1]\, B => 
        \asize_reg[0]_net_1\, C => \RDATA_reg[17]_net_1\, Y => 
        m30_1_1_2);
    
    \WDATA_reg[0]\ : SLE
      port map(D => \WDATA_mux[0]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[0]_net_1\);
    
    \WSTRB_mux_3_0[3]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \WSTRB_reg[3]_net_1\, B => 
        \WSTRB_mux_3_0_a3_0_0[3]_net_1\, C => N_3149_2, D => 
        N_3141, Y => \WSTRB_mux[3]\);
    
    \WDATA_mux_3_0[13]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[13]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[13]_net_1\, Y => \WDATA_mux[13]\);
    
    raddr_reg_9_2_axb_20_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(21), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(21), Y => 
        \raddr_reg_9_2_axb_20_1\);
    
    \axi_state[8]\ : SLE
      port map(D => \axi_state_ns[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_ARREADY\);
    
    raddr_reg_9_2_axb_15_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(16), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(16), Y => 
        \raddr_reg_9_2_axb_15_1\);
    
    \RDATA_reg_RNO[55]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[55]_net_1\, D => 
        \sdr_dataout_reg[7]_net_1\, Y => N_193_mux_i);
    
    \RDATA_reg_RNI17GJ1[16]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[16]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[0]\, C => N_3141, D => 
        N_3167_i, Y => N_72_mux_i);
    
    \raddr_reg[1]\ : SLE
      port map(D => \raddr_reg_9[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[1]_net_1\);
    
    \asize[1]\ : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARSIZE(1), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWSIZE(1), Y => \asize[1]_net_1\);
    
    \WDATA_mux_31[18]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(50), B => 
        COREAXI_0_AXImslave16_WDATA(18), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[18]_net_1\);
    
    \sdr_datain_2[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[11]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[11]_net_1\);
    
    \WDATA_reg[18]\ : SLE
      port map(D => \WDATA_mux[18]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[18]_net_1\);
    
    \WDATA_mux_15_3[15]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(15), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[15]_net_1\);
    
    \raddr_reg_RNIV17V7[4]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[4]_net_1\, C => 
        \raddr_reg_9_2_axb_4_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_3, S => N_753, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_4);
    
    \raddr_reg_9[15]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_764, Y => \raddr_reg_9[15]_net_1\);
    
    \sdr_datain_reg[2]\ : SLE
      port map(D => \sdr_datain[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(2));
    
    \raddr_reg[15]\ : SLE
      port map(D => \raddr_reg_9[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[15]_net_1\);
    
    \raddr_reg[0]\ : SLE
      port map(D => \raddr_reg_9[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[0]_net_1\);
    
    \sdr_datain_reg_RNO[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[3]_net_1\, C => \sdr_datain_1[3]_net_1\, Y
         => \sdr_datain[3]\);
    
    \sdr_dataout_reg[8]\ : SLE
      port map(D => DQ_in(8), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[8]_net_1\);
    
    \WDATA_reg[52]\ : SLE
      port map(D => \WDATA_mux[52]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[52]_net_1\);
    
    \sdr_datain_0[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[17]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[1]_net_1\);
    
    \RDATA_reg[0]\ : SLE
      port map(D => N_170_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[0]\);
    
    \B_SIZE_reg_RNIESI41[0]\ : CFG4
      generic map(INIT => x"EB7D")

      port map(A => \B_SIZE_reg[0]_net_1\, B => 
        \B_SIZE_reg[1]_net_1\, C => \sdr_count[1]_net_1\, D => 
        \sdr_count[0]_net_1\, Y => un2_sdr_count_NE_0);
    
    \RDATA_reg[20]\ : SLE
      port map(D => \sdr_dataout_reg[4]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[20]_net_1\);
    
    \raddr_reg[2]\ : SLE
      port map(D => \raddr_reg_9[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[2]_net_1\);
    
    \raddr_reg[19]\ : SLE
      port map(D => \raddr_reg_9[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[19]_net_1\);
    
    \WDATA_mux_3_0_RNO[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[1]_net_1\, C => \WDATA_mux_8_1[1]_net_1\, 
        Y => \WDATA_mux_8[1]\);
    
    \WDATA_mux_31[21]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(53), B => 
        COREAXI_0_AXImslave16_WDATA(21), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[21]_net_1\);
    
    \WDATA_reg[62]\ : SLE
      port map(D => \WDATA_mux[62]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[62]_net_1\);
    
    \WDATA_mux_3_0[7]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[7]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[7]_net_1\, Y => \WDATA_mux[7]\);
    
    \RDATA_reg[12]\ : SLE
      port map(D => N_182_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[12]\);
    
    \WDATA_mux_3_0_RNO[12]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[12]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[12]_net_1\, Y => \WDATA_mux_15[12]\);
    
    un1_sdr_count_0_sqmuxa_0 : CFG4
      generic map(INIT => x"FCF8")

      port map(A => \axi_state[3]_net_1\, B => W_VALID, C => 
        N_358, D => \axi_state[0]_net_1\, Y => 
        un1_sdr_count_0_sqmuxa);
    
    WE_N : SLE
      port map(D => WE_N_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => WE_N_c);
    
    \RDATA_reg_RNIVQGN1[56]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[56]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_1_i_1);
    
    \raddr_reg_RNITCM6M[15]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[15]_net_1\, C => 
        \raddr_reg_9_2_axb_15_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_14, S => N_764, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_15);
    
    \RDATA_reg[43]\ : SLE
      port map(D => \sdr_dataout_reg[11]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_reg_0);
    
    \WDATA_mux_15_1[9]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[9]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(25), D
         => COREAXI_0_AXImslave16_WDATA(41), Y => 
        \WDATA_mux_15_1[9]_net_1\);
    
    \sdr_datain_0[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[31]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[15]_net_1\);
    
    \asize_reg_RNIEK505[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_8\, C => i22_mux_1_i_1_0, 
        D => i22_mux_1_i_1, Y => i22_mux_1_i);
    
    \sdr_datain_reg[10]\ : SLE
      port map(D => \sdr_datain[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(10));
    
    \raddr_reg_9[21]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_770, Y => \raddr_reg_9[21]_net_1\);
    
    \WDATA_mux_3_0_RNO[15]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[15]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[15]_net_1\, Y => \WDATA_mux_15[15]\);
    
    \axi_state_ns_i_0[4]\ : CFG4
      generic map(INIT => x"A0EC")

      port map(A => COREAXI_0_AXImslave16_WVALID, B => 
        \COREAXI_0_AXImslave16_AWREADY\, C => 
        \axi_state[5]_net_1\, D => COREAXI_0_AXImslave16_AWVALID, 
        Y => \axi_state_ns_i_0[4]_net_1\);
    
    \RDATA_reg[3]\ : SLE
      port map(D => N_173_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[3]\);
    
    \RDATA_reg_RNIVNDN1[29]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[29]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_1_i_1_0);
    
    \raddr_reg_9[12]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_761, Y => \raddr_reg_9[12]_net_1\);
    
    \WDATA_mux_3_0_a2_0[15]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \asize_reg[0]_net_1\, B => 
        \asize_reg[1]_net_1\, C => COREAXI_0_AXImslave16_WSTRB(1), 
        D => COREAXI_0_AXImslave16_WSTRB(5), Y => N_3236);
    
    \WDATA_mux_3_0[10]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[10]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[10]_net_1\, Y => \WDATA_mux[10]\);
    
    \RDATA_reg_RNO[4]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[4]\, D => 
        \sdr_dataout_reg[4]_net_1\, Y => N_174_mux_i);
    
    \RDATA_reg[27]\ : SLE
      port map(D => \sdr_dataout_reg[11]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[27]_net_1\);
    
    \sdr_dataout_reg[6]\ : SLE
      port map(D => DQ_in(6), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[6]_net_1\);
    
    \WDATA_mux_8_1[5]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[5]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(37), D
         => COREAXI_0_AXImslave16_WDATA(21), Y => 
        \WDATA_mux_8_1[5]_net_1\);
    
    \sdr_count_RNI201B[3]\ : CFG4
      generic map(INIT => x"EEEF")

      port map(A => \sdr_count[2]_net_1\, B => 
        \sdr_count[3]_net_1\, C => \sdr_count[1]_net_1\, D => 
        \sdr_count[0]_net_1\, Y => \sdr_count_RNI201B[3]_net_1\);
    
    \WDATA_reg_RNO[41]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(41), 
        Y => \WDATA_mux[41]\);
    
    \WDATA_mux_8_3[1]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(1), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[1]_net_1\);
    
    \sdr_dataout_reg[2]\ : SLE
      port map(D => DQ_in(2), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[2]_net_1\);
    
    \axi_state[3]\ : SLE
      port map(D => N_311_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[3]_net_1\);
    
    \sdr_datain_reg[1]\ : SLE
      port map(D => \sdr_datain[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(1));
    
    \axi_state[9]\ : SLE
      port map(D => \axi_state_ns[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[9]_net_1\);
    
    \WDATA_reg[50]\ : SLE
      port map(D => \WDATA_mux[50]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[50]_net_1\);
    
    \RDATA_reg_RNIUMDN1[28]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[28]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_i_1_0);
    
    \raddr_reg_RNID9LSC[8]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[8]_net_1\, C => 
        \raddr_reg_9_2_axb_8_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_7, S => N_757, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_8);
    
    \sdr_datain_2[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[3]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[3]_net_1\);
    
    \sdr_datain_0[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[28]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[12]_net_1\);
    
    \RDATA_reg_RNO[54]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[54]_net_1\, D => 
        \sdr_dataout_reg[6]_net_1\, Y => N_192_mux_i);
    
    raddr_reg_9_2_axb_13_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(14), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(14), Y => 
        \raddr_reg_9_2_axb_13_1\);
    
    \axi_state_ns_0[5]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_BVALID, B => 
        N_3309, C => \COREAXI_0_AXImslave16_BVALID\, Y => 
        \axi_state_ns[5]\);
    
    \RDATA_reg[24]\ : SLE
      port map(D => \sdr_dataout_reg[8]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[24]_net_1\);
    
    \B_SIZE_reg[2]\ : SLE
      port map(D => b_size4, CLK => SDRCLK_c, EN => N_295_i, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \B_SIZE_reg[2]_net_1\);
    
    \RDATA_reg_RNO[12]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[12]\, D => 
        \sdr_dataout_reg[12]_net_1\, Y => N_182_mux_i);
    
    \sdr_dataout_reg[4]\ : SLE
      port map(D => DQ_in(4), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[4]_net_1\);
    
    \asize_reg_RNIRE215[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_13\, C => i17_mux_1_i_1_0, 
        D => i17_mux_1_i_1, Y => i17_mux_1_i);
    
    \WDATA_reg[60]\ : SLE
      port map(D => \WDATA_mux[60]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[60]_net_1\);
    
    \sdr_dataout_reg[15]\ : SLE
      port map(D => DQ_in(15), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[15]_net_1\);
    
    \sdr_datain_1[6]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[6]_net_1\, C => \WDATA_reg[54]_net_1\, D
         => \WDATA_reg[38]_net_1\, Y => \sdr_datain_1[6]_net_1\);
    
    \RDATA_reg_RNICRFQ1[38]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[6]\, B => 
        \RDATA_reg[38]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3098_i);
    
    \RDATA_reg_RNIMEDN1[20]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[20]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_5_i_1_0);
    
    \RDATA_reg[10]\ : SLE
      port map(D => N_180_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[10]\);
    
    \raddr_reg_RNI780OG[11]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[11]_net_1\, C => 
        \raddr_reg_9_2_axb_11_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_10, S => N_760, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_11);
    
    \un1_B_SIZE_reg_0_a2_RNISOQQ1[2]\ : ARI1
      generic map(INIT => x"5758A")

      port map(A => \raddr_reg_RNIOTA71[0]_net_1\, B => 
        \un1_B_SIZE_reg_0_a2[2]_net_1\, C => N_335_i, D => 
        \axi_state[9]_net_1\, FCI => GND_net_1, S => OPEN, Y => 
        \un1_B_SIZE_reg_0_a2_RNISOQQ1_Y[2]\, FCO => 
        raddr_reg_9_2_cry_0);
    
    raddr_reg_9_2_axb_17_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(18), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(18), Y => 
        \raddr_reg_9_2_axb_17_1\);
    
    \WDATA_mux_15_0[11]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(59), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[11]_net_1\);
    
    \raddr_reg_9[5]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_754, Y => \raddr_reg_9[5]_net_1\);
    
    \WSTRB_reg[6]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(6), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[6]_net_1\);
    
    \RDATA_reg_RNO[60]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[60]_net_1\, D => 
        \sdr_dataout_reg[12]_net_1\, Y => N_198_mux_i);
    
    \RDATA_reg_RNI6APC1[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[10]\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_10);
    
    \WDATA_mux_3_0_0[13]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(13), B => 
        COREAXI_0_AXImslave16_WDATA(45), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[13]_net_1\);
    
    \raddr_reg_9[16]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_765, Y => \raddr_reg_9[16]_net_1\);
    
    \sdr_dataout_reg[0]\ : SLE
      port map(D => DQ_in(0), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[0]_net_1\);
    
    \RDATA_reg_RNI4JFQ1[34]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[2]\, B => 
        \RDATA_reg[34]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_34);
    
    \RDATA_reg_RNIHQQQ[49]\ : CFG4
      generic map(INIT => x"7D41")

      port map(A => \RDATA_reg[49]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        m30_1_1_2, Y => i58_mux_2);
    
    \SA[9]\ : SLE
      port map(D => \SA_i[9]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(9));
    
    \sdr_datain_3[11]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[11]_net_1\, C => \WDATA_reg[11]_net_1\, Y
         => \sdr_datain_3[11]_net_1\);
    
    un61_axi_state_i_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \R_VALID\, B => W_VALID, Y => N_388);
    
    \WDATA_reg_RNO[52]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(52), 
        Y => \WDATA_mux[52]\);
    
    \WDATA_reg[57]\ : SLE
      port map(D => \WDATA_mux[57]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[57]_net_1\);
    
    \WDATA_reg[21]\ : SLE
      port map(D => \WDATA_mux[21]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[21]_net_1\);
    
    \sdr_datain_1[15]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[15]_net_1\, C => \WDATA_reg[63]_net_1\, D
         => \WDATA_reg[47]_net_1\, Y => \sdr_datain_1[15]_net_1\);
    
    \asize_reg_RNIUG115[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_11\, C => i22_mux_0_i_1_0, 
        D => i22_mux_0_i_1, Y => i22_mux_0_i);
    
    \WDATA_reg[43]\ : SLE
      port map(D => \WDATA_mux[43]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[43]_net_1\);
    
    \WDATA_mux_3_0_m4[7]\ : CFG3
      generic map(INIT => x"AD")

      port map(A => \asize_reg[1]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(0), C => \asize_reg[0]_net_1\, 
        Y => N_3240);
    
    \RDATA_reg[33]\ : SLE
      port map(D => \sdr_dataout_reg[1]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[33]_net_1\);
    
    \RDATA_reg_RNI9PGQ1[41]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[9]\, B => 
        \RDATA_reg[41]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_41);
    
    \WDATA_reg_RNO[63]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(63), 
        Y => \WDATA_mux[63]\);
    
    \WDATA_mux_3_0_RNO[7]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[7]_net_1\, C => \WDATA_mux_8_1[7]_net_1\, 
        Y => \WDATA_mux_8[7]\);
    
    \axi_state_ns_0[7]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => \axi_state_0\, B => N_23, C => 
        \axi_state_ns_0_0[7]_net_1\, D => \N_3297\, Y => 
        \axi_state_ns[7]\);
    
    \RDATA_reg[17]\ : SLE
      port map(D => N_3070_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[17]_net_1\);
    
    \WDATA_mux_3_0_0[5]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(5), B => 
        COREAXI_0_AXImslave16_WDATA(37), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[5]_net_1\);
    
    \asize_reg[0]\ : SLE
      port map(D => \asize_reg_134\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \asize_reg[0]_net_1\);
    
    \sdr_datain_2[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[10]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[10]_net_1\);
    
    \WDATA_reg[54]\ : SLE
      port map(D => \WDATA_mux[54]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[54]_net_1\);
    
    \SA[4]\ : SLE
      port map(D => \SA_i[4]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(4));
    
    \WDATA_reg_RNO[45]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(45), 
        Y => \WDATA_mux[45]\);
    
    \sdr_datain_1[7]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[7]_net_1\, C => \WDATA_reg[55]_net_1\, D
         => \WDATA_reg[39]_net_1\, Y => \sdr_datain_1[7]_net_1\);
    
    raddr_reg_9_2_axb_18_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(19), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(19), Y => 
        \raddr_reg_9_2_axb_18_1\);
    
    \axi_state_RNO[3]\ : CFG4
      generic map(INIT => x"A8FC")

      port map(A => \axi_state[5]_net_1\, B => \WREADY_SI16\, C
         => \axi_state[3]_net_1\, D => RW_ACK, Y => N_311_i);
    
    \sdr_datain_1[12]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[12]_net_1\, C => \WDATA_reg[60]_net_1\, D
         => \WDATA_reg[44]_net_1\, Y => \sdr_datain_1[12]_net_1\);
    
    \raddr_reg_9[13]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_762, Y => \raddr_reg_9[13]_net_1\);
    
    \raddr_reg_9[11]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_760, Y => \raddr_reg_9[11]_net_1\);
    
    \WDATA_mux_3_0_0[0]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(0), B => 
        COREAXI_0_AXImslave16_WDATA(32), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[0]_net_1\);
    
    \WDATA_mux_15_1[13]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[13]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(29), D
         => COREAXI_0_AXImslave16_WDATA(45), Y => 
        \WDATA_mux_15_1[13]_net_1\);
    
    \RDATA_reg[14]\ : SLE
      port map(D => N_184_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA_3\);
    
    \asize_reg[1]\ : SLE
      port map(D => \asize_reg_135\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \asize_reg[1]_net_1\);
    
    \WDATA_mux_15_3[8]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(8), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[8]_net_1\);
    
    \WDATA_mux_3_0_RNO[10]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[10]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[10]_net_1\, Y => \WDATA_mux_15[10]\);
    
    \WDATA_mux_3_0_RNO[14]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[14]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[14]_net_1\, Y => \WDATA_mux_15[14]\);
    
    \sdr_datain_2[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[13]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[13]_net_1\);
    
    \sdr_datain_1[4]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[4]_net_1\, C => \WDATA_reg[52]_net_1\, D
         => \WDATA_reg[36]_net_1\, Y => \sdr_datain_1[4]_net_1\);
    
    \WDATA_reg[13]\ : SLE
      port map(D => \WDATA_mux[13]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[13]_net_1\);
    
    \WDATA_mux_3[22]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(22), C => 
        \WDATA_mux_31[22]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[22]\);
    
    \un7_1.N_3272_i\ : CFG4
      generic map(INIT => x"0A09")

      port map(A => \axi_count[2]_net_1\, B => 
        \axi_count[1]_net_1\, C => N_3293, D => N_3289, Y => 
        N_3272_i);
    
    \WDATA_reg_RNO[33]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(33), 
        Y => \WDATA_mux[33]\);
    
    \WDATA_reg[38]\ : SLE
      port map(D => \WDATA_mux[38]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[38]_net_1\);
    
    \RDATA_reg_RNIL8DK1[27]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[27]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_0\, C => N_3141, D => 
        N_3167_i, Y => N_76_mux_i);
    
    \sdr_count[0]\ : SLE
      port map(D => N_3280_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_count[0]_net_1\);
    
    \axi_state_ns[2]\ : CFG4
      generic map(INIT => x"C202")

      port map(A => \COREAXI_0_AXImslave16_AWREADY\, B => 
        COREAXI_0_AXImslave16_AWVALID, C => \axi_state[9]_net_1\, 
        D => un5_axi_rvalid_i_0, Y => \axi_state_ns[2]_net_1\);
    
    \axi_count[0]\ : SLE
      port map(D => N_3276_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_count[0]_net_1\);
    
    \RDATA_reg[52]\ : SLE
      port map(D => N_190_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[52]_net_1\);
    
    \sdr_datain_1[1]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[1]_net_1\, C => \WDATA_reg[49]_net_1\, D
         => \WDATA_reg[33]_net_1\, Y => \sdr_datain_1[1]_net_1\);
    
    \WDATA_mux_3[23]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(23), C => 
        \WDATA_mux_31[23]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[23]\);
    
    \WDATA_mux_15_0[10]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(58), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[10]_net_1\);
    
    \WSTRB_reg_RNIA8EL[6]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \WSTRB_reg[7]_net_1\, B => 
        \WSTRB_reg[6]_net_1\, C => \WSTRB_reg[5]_net_1\, D => 
        \WSTRB_reg[4]_net_1\, Y => WSTRB_mux_8_sn_m3_i_a3_1);
    
    \WDATA_mux_3_0_0[3]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(3), B => 
        COREAXI_0_AXImslave16_WDATA(35), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[3]_net_1\);
    
    \SA[7]\ : SLE
      port map(D => \SA_i[7]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(7));
    
    \raddr_reg_RNIQ5CIN[16]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[16]_net_1\, C => 
        \raddr_reg_9_2_axb_16_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_15, S => N_765, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_16);
    
    \WSTRB_reg[7]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(7), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[7]_net_1\);
    
    \RDATA_reg[26]\ : SLE
      port map(D => \sdr_dataout_reg[10]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[26]_net_1\);
    
    \axi_count[2]\ : SLE
      port map(D => N_3272_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_count[2]_net_1\);
    
    asize_reg_0_sqmuxa_i : CFG3
      generic map(INIT => x"A8")

      port map(A => \axi_state[9]_net_1\, B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWVALID, Y => N_295_i);
    
    \axi_state_ns[1]\ : CFG4
      generic map(INIT => x"02CE")

      port map(A => \COREAXI_0_AXImslave16_ARREADY\, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => un5_axi_rvalid_i_0, Y => \axi_state_ns[1]_net_1\);
    
    \sdr_datain_2[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[5]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[5]_net_1\);
    
    \RDATA_reg_RNI39GJ1[17]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[17]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[1]\, C => N_3141, D => 
        N_3167_i, Y => N_71_mux_i);
    
    \WDATA_mux_3_0_0[8]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(8), B => 
        COREAXI_0_AXImslave16_WDATA(40), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[8]_net_1\);
    
    \sdr_dataout_reg[10]\ : SLE
      port map(D => DQ_in(10), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[10]_net_1\);
    
    \sdr_datain_2[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[7]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[7]_net_1\);
    
    \WDATA_mux_3_0[5]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[5]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[5]_net_1\, Y => \WDATA_mux[5]\);
    
    \sdr_datain_reg[15]\ : SLE
      port map(D => \sdr_datain[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(15));
    
    \RDATA_reg_RNI5BGJ1[18]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[18]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[2]\, C => N_3141, D => 
        N_3167_i, Y => N_70_mux_i);
    
    \SA[8]\ : SLE
      port map(D => \SA_i[8]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(8));
    
    \WDATA_mux_8_0[7]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(55), B => 
        COREAXI_0_AXImslave16_WSTRB(6), C => 
        COREAXI_0_AXImslave16_WSTRB(4), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[7]_net_1\);
    
    \RDATA_reg_RNIMICR1[44]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[12]\, B => 
        \RDATA_reg[44]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3092_i);
    
    \RDATA_reg_RNO[18]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[18]_net_1\, D => 
        \sdr_dataout_reg[2]_net_1\, Y => N_3071_i);
    
    \raddr_reg_9_2_1_1[0]\ : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(1), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(1), Y => 
        \raddr_reg_9_2_1_1[0]_net_1\);
    
    \WDATA_mux_3_0[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(62), B => 
        COREAXI_0_AXImslave16_WDATA(30), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[30]\);
    
    \WDATA_reg_RNO[39]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(39), 
        Y => \WDATA_mux[39]\);
    
    \WDATA_mux_15_3[11]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(11), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[11]_net_1\);
    
    raddr_reg_9_2_axb_9_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(10), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(10), Y => 
        \raddr_reg_9_2_axb_9_1\);
    
    \WDATA_reg_RNO[44]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(44), 
        Y => \WDATA_mux[44]\);
    
    \sdr_datain_0[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[27]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[11]_net_1\);
    
    \WDATA_reg[56]\ : SLE
      port map(D => \WDATA_mux[56]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[56]_net_1\);
    
    \RDATA_reg[50]\ : SLE
      port map(D => N_188_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[50]_net_1\);
    
    \WDATA_reg_RNO[58]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(58), 
        Y => \WDATA_mux[58]\);
    
    \sdr_datain_3[10]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[10]_net_1\, C => \WDATA_reg[10]_net_1\, Y
         => \sdr_datain_3[10]_net_1\);
    
    \un1_B_SIZE_reg_0_a2_RNIQGGG5[0]\ : ARI1
      generic map(INIT => x"5758A")

      port map(A => \raddr_reg_RNIU3B71[2]_net_1\, B => 
        \un1_B_SIZE_reg_0_a2[0]_net_1\, C => N_335_i, D => 
        \axi_state[9]_net_1\, FCI => raddr_reg_9_2_cry_1, S => 
        N_751, Y => OPEN, FCO => raddr_reg_9_2_cry_2);
    
    \WDATA_mux_15_1[14]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[14]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(30), D
         => COREAXI_0_AXImslave16_WDATA(46), Y => 
        \WDATA_mux_15_1[14]_net_1\);
    
    \RDATA_reg[2]\ : SLE
      port map(D => N_172_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[2]\);
    
    \sdr_datain_reg_RNO[10]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[10]_net_1\, C => \sdr_datain_1[10]_net_1\, 
        Y => \sdr_datain[10]\);
    
    \sdr_count_RNO[0]\ : CFG4
      generic map(INIT => x"0014")

      port map(A => N_3281, B => un1_sdr_count_0_sqmuxa, C => 
        \sdr_count[0]_net_1\, D => N_3293, Y => N_3280_i);
    
    \WSTRB_mux_3_0_m3[1]\ : CFG4
      generic map(INIT => x"AAAC")

      port map(A => \WSTRB_reg[1]_net_1\, B => 
        \WSTRB_mux_8_m1[1]_net_1\, C => N_3141, D => N_26, Y => 
        N_3144);
    
    \RDATA_reg[16]\ : SLE
      port map(D => N_3069_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[16]_net_1\);
    
    \raddr_reg_RNIHIFLR[19]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[19]_net_1\, C => 
        \raddr_reg_9_2_axb_19_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_18, S => N_768, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_19);
    
    \WSTRB_mux_3_0_o3[3]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \asize_reg[1]_net_1\, B => 
        \asize_reg[0]_net_1\, Y => N_3141);
    
    \WDATA_mux_15_1[8]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[8]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(24), D
         => COREAXI_0_AXImslave16_WDATA(40), Y => 
        \WDATA_mux_15_1[8]_net_1\);
    
    \axi_state[5]\ : SLE
      port map(D => N_308_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[5]_net_1\);
    
    \raddr_reg[16]\ : SLE
      port map(D => \raddr_reg_9[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[16]_net_1\);
    
    \RDATA_reg_RNO[29]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[29]_net_1\, D => 
        \sdr_dataout_reg[13]_net_1\, Y => N_3072_i);
    
    \RDATA_reg_RNO[10]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[10]\, D => 
        \sdr_dataout_reg[10]_net_1\, Y => N_180_mux_i);
    
    \SA[6]\ : SLE
      port map(D => \SA_i[6]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(6));
    
    \xhdl21.b_size3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \asize[1]_net_1\, B => \asize[0]_net_1\, Y
         => b_size3);
    
    \sdr_datain_3[13]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[13]_net_1\, C => \WDATA_reg[13]_net_1\, Y
         => \sdr_datain_3[13]_net_1\);
    
    un3_r_req_0_0 : CFG3
      generic map(INIT => x"EA")

      port map(A => \axi_state[2]_net_1\, B => \axi_state_0\, C
         => N_23, Y => \un3_r_req_0_0\);
    
    \sdr_datain_reg_RNO[7]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[7]_net_1\, C => \sdr_datain_1[7]_net_1\, Y
         => \sdr_datain[7]\);
    
    \sdr_datain_3[7]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[7]_net_1\, C => \WDATA_reg[7]_net_1\, Y => 
        \sdr_datain_3[7]_net_1\);
    
    \WDATA_mux_3_0_0[9]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(9), B => 
        COREAXI_0_AXImslave16_WDATA(41), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[9]_net_1\);
    
    un1_rvalid_xhdl1_i_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \axi_count[2]_net_1\, B => 
        \axi_count[3]_net_1\, C => \axi_count[1]_net_1\, D => 
        \axi_count[0]_net_1\, Y => \N_389\);
    
    \WDATA_mux_3_0_RNO[11]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[11]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[11]_net_1\, Y => \WDATA_mux_15[11]\);
    
    \RDATA_reg[57]\ : SLE
      port map(D => N_195_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[57]_net_1\);
    
    \RDATA_reg[29]\ : SLE
      port map(D => N_3072_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[29]_net_1\);
    
    \RDATA_reg_RNIUPGN1[55]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[55]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_2_i_1);
    
    \WDATA_mux_3_0[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(58), B => 
        COREAXI_0_AXImslave16_WDATA(26), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[26]\);
    
    \sdr_datain_2[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[14]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[14]_net_1\);
    
    \raddr_reg_9[4]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_753, Y => \raddr_reg_9[4]_net_1\);
    
    \WDATA_reg_RNO[50]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(50), 
        Y => \WDATA_mux[50]\);
    
    \RDATA_reg_RNO[49]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[49]_net_1\, D => 
        \sdr_dataout_reg[1]_net_1\, Y => N_187_mux_i);
    
    \sdr_datain_reg[12]\ : SLE
      port map(D => \sdr_datain[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(12));
    
    \RDATA_reg[42]\ : SLE
      port map(D => \sdr_dataout_reg[10]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[42]_net_1\);
    
    \sdr_datain_reg[0]\ : SLE
      port map(D => \sdr_datain[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(0));
    
    \RDATA_reg_RNO[57]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[57]_net_1\, D => 
        \sdr_dataout_reg[9]_net_1\, Y => N_195_mux_i);
    
    \WSTRB_reg[5]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(5), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[5]_net_1\);
    
    \WDATA_mux_3_0[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(57), B => 
        COREAXI_0_AXImslave16_WDATA(25), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[25]\);
    
    \RDATA_reg_RNIBLRQ[50]\ : CFG4
      generic map(INIT => x"7D41")

      port map(A => \RDATA_reg[50]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        m23_1_2, Y => i58_mux_1);
    
    \RDATA_reg[54]\ : SLE
      port map(D => N_192_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[54]_net_1\);
    
    \B_SIZE_reg[0]\ : SLE
      port map(D => \asize[1]_net_1\, CLK => SDRCLK_c, EN => 
        N_295_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \B_SIZE_reg[0]_net_1\);
    
    \WDATA_mux_8_1[7]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[7]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(39), D
         => COREAXI_0_AXImslave16_WDATA(23), Y => 
        \WDATA_mux_8_1[7]_net_1\);
    
    \WDATA_mux_15_1[15]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[15]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(31), D
         => COREAXI_0_AXImslave16_WDATA(47), Y => 
        \WDATA_mux_15_1[15]_net_1\);
    
    R_VALID_reg : SLE
      port map(D => R_VALID_i, CLK => SDRCLK_c, EN => MSS_READY, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \R_VALID_reg\);
    
    \sdr_datain_1[11]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[11]_net_1\, C => \WDATA_reg[59]_net_1\, D
         => \WDATA_reg[43]_net_1\, Y => \sdr_datain_1[11]_net_1\);
    
    \sdr_datain_0[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[19]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[3]_net_1\);
    
    \RDATA_reg_RNO[3]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[3]\, D => 
        \sdr_dataout_reg[3]_net_1\, Y => N_173_mux_i);
    
    \WDATA_mux_15_3[10]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(10), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[10]_net_1\);
    
    \raddr_reg[6]\ : SLE
      port map(D => \raddr_reg_9[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[6]_net_1\);
    
    R_VALID : SLE
      port map(D => \R_VALID_reg\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \R_VALID\);
    
    \WDATA_mux_3_0_0[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(11), B => 
        COREAXI_0_AXImslave16_WDATA(43), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[11]_net_1\);
    
    \sdr_datain_reg[13]\ : SLE
      port map(D => \sdr_datain[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(13));
    
    \WDATA_reg_RNO[61]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(61), 
        Y => \WDATA_mux[61]\);
    
    \RDATA_regce[32]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \sdr_count[1]_net_1\, B => \R_VALID\, C => 
        \sdr_count[0]_net_1\, Y => \RDATA_regce[32]_net_1\);
    
    \RDATA_reg_RNIOHEN1[31]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[31]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_i_1_0);
    
    \sdr_count_RNO[3]\ : CFG4
      generic map(INIT => x"0A06")

      port map(A => \sdr_count[3]_net_1\, B => 
        \sdr_count[2]_net_1\, C => N_3299, D => N_3288, Y => 
        N_3277_i);
    
    \raddr_reg_RNIGE0DU[21]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[21]_net_1\, C => 
        \raddr_reg_9_2_axb_21_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_20, S => N_770, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_21);
    
    \WDATA_mux_3_0[8]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[8]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[8]_net_1\, Y => \WDATA_mux[8]\);
    
    \asize_reg_RNI8C305[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_0\, C => i17_mux_2_i_1_0, 
        D => i17_mux_2_i_1, Y => i17_mux_2_i);
    
    \WSTRB_reg_RNIU7381[0]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => \un7_wstrb_reg_i_a3\, B => 
        WSTRB_mux_8_sn_m3_i_a3_1, C => \WSTRB_reg[1]_net_1\, D
         => \WSTRB_reg[0]_net_1\, Y => N_26);
    
    \WDATA_reg[59]\ : SLE
      port map(D => \WDATA_mux[59]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[59]_net_1\);
    
    \WDATA_reg[2]\ : SLE
      port map(D => \WDATA_mux[2]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[2]_net_1\);
    
    \sdr_datain_2[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[1]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[1]_net_1\);
    
    \WDATA_reg[33]\ : SLE
      port map(D => \WDATA_mux[33]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[33]_net_1\);
    
    raddr_reg_9_2_axb_5_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(6), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(6), Y => 
        \raddr_reg_9_2_axb_5_1\);
    
    raddr_reg_9_2_axb_10_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(11), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(11), Y => 
        \raddr_reg_9_2_axb_10_1\);
    
    \RDATA_reg_RNO[16]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[16]_net_1\, D => 
        \sdr_dataout_reg[0]_net_1\, Y => N_3069_i);
    
    \axi_state_ns_0_a2[0]\ : CFG3
      generic map(INIT => x"40")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => un5_axi_rvalid_i_0, Y => 
        N_3313);
    
    \WDATA_reg[28]\ : SLE
      port map(D => \WDATA_mux[28]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[28]_net_1\);
    
    \RDATA_reg[19]\ : SLE
      port map(D => \sdr_dataout_reg[3]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[19]_net_1\);
    
    \RDATA_reg[61]\ : SLE
      port map(D => N_199_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[61]_net_1\);
    
    CKE : SLE
      port map(D => CKE_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => CKE_c);
    
    \RDATA_reg_RNISNGN1[53]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[53]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_4_i_1);
    
    \RDATA_reg[25]\ : SLE
      port map(D => \sdr_dataout_reg[9]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[25]_net_1\);
    
    \RDATA_reg_RNITKTB1[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[8]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_8\);
    
    \DQM[1]\ : SLE
      port map(D => \DQM_i_3[1]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        DQM_c(1));
    
    \RDATA_reg[40]\ : SLE
      port map(D => \sdr_dataout_reg[8]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[40]_net_1\);
    
    \WDATA_mux_3_0_RNO[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[5]_net_1\, C => \WDATA_mux_8_1[5]_net_1\, 
        Y => \WDATA_mux_8[5]\);
    
    \B_SIZE_reg[1]\ : SLE
      port map(D => b_size3, CLK => SDRCLK_c, EN => N_295_i, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \B_SIZE_reg[1]_net_1\);
    
    \sdr_datain_3[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[4]_net_1\, C => \WDATA_reg[4]_net_1\, Y => 
        \sdr_datain_3[4]_net_1\);
    
    \sdr_datain_1[0]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[0]_net_1\, C => \WDATA_reg[48]_net_1\, D
         => \WDATA_reg[32]_net_1\, Y => \sdr_datain_1[0]_net_1\);
    
    \WDATA_reg_RNO[56]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(56), 
        Y => \WDATA_mux[56]\);
    
    \WDATA_mux_3_0[28]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(60), B => 
        COREAXI_0_AXImslave16_WDATA(28), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[28]\);
    
    \WDATA_reg[42]\ : SLE
      port map(D => \WDATA_mux[42]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[42]_net_1\);
    
    \raddr_reg_9[3]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_752, Y => \raddr_reg_9[3]_net_1\);
    
    \WSTRB_mux_3_0_a3_0_2[2]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \WSTRB_reg[0]_net_1\, B => 
        \WSTRB_reg[1]_net_1\, C => \asize_reg[0]_net_1\, D => 
        \asize_reg[1]_net_1\, Y => N_3149_2);
    
    \RDATA_reg_RNIEC4D[26]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \COREAXI_0_AXImslave16_RDATA[10]\, B => 
        \asize_reg[0]_net_1\, C => \RDATA_reg[26]_net_1\, Y => 
        m9_1_1_2);
    
    \un7_1.SUM_i_o2_2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \axi_count[1]_net_1\, B => 
        \axi_count[2]_net_1\, Y => N_3286);
    
    \RDATA_reg_RNI7NGQ1[40]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[8]\, B => 
        \RDATA_reg[40]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3094_i);
    
    \RDATA_reg[32]\ : SLE
      port map(D => \sdr_dataout_reg[0]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[32]_net_1\);
    
    \WDATA_reg[4]\ : SLE
      port map(D => \WDATA_mux[4]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[4]_net_1\);
    
    \sdr_datain_0[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[26]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[10]_net_1\);
    
    \DQM_mux_ns_1[1]\ : CFG4
      generic map(INIT => x"5702")

      port map(A => \sdr_count[1]_net_1\, B => 
        \DQM_mux_ns_1_1[1]_net_1\, C => \N_74\, D => 
        \WSTRB_mux[3]\, Y => \DQM_mux_ns_1[1]_net_1\);
    
    \axi_state[1]\ : SLE
      port map(D => \axi_state_ns[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_state[1]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \RDATA_reg_RNI9DPC1[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[13]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_13\);
    
    \WDATA_mux_3_0_0[1]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(1), B => 
        COREAXI_0_AXImslave16_WDATA(33), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[1]_net_1\);
    
    \axi_state_RNO[5]\ : CFG4
      generic map(INIT => x"000D")

      port map(A => \N_389\, B => \COREAXI_0_AXImslave16_AWREADY\, 
        C => N_368, D => \axi_state_ns_i_0[4]_net_1\, Y => 
        N_308_i);
    
    \sdr_datain_1[9]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[9]_net_1\, C => \WDATA_reg[57]_net_1\, D
         => \WDATA_reg[41]_net_1\, Y => \sdr_datain_1[9]_net_1\);
    
    \WDATA_mux_15_0[12]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(60), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[12]_net_1\);
    
    \WDATA_mux_8_1[0]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => WDATA_mux_8_sm0, B => 
        \WDATA_mux_8_0[0]_net_1\, C => 
        COREAXI_0_AXImslave16_WDATA(16), D => 
        COREAXI_0_AXImslave16_WDATA(32), Y => 
        \WDATA_mux_8_1[0]_net_1\);
    
    \RDATA_reg[47]\ : SLE
      port map(D => \sdr_dataout_reg[15]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[47]_net_1\);
    
    \raddr_reg_9[8]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_757, Y => \raddr_reg_9[8]_net_1\);
    
    \sdr_datain_3[14]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[14]_net_1\, C => \WDATA_reg[14]_net_1\, Y
         => \sdr_datain_3[14]_net_1\);
    
    \WDATA_mux_3_0_0[7]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(7), B => 
        COREAXI_0_AXImslave16_WDATA(39), C => N_3240, D => N_3268, 
        Y => \WDATA_mux_3_0_0[7]_net_1\);
    
    \RDATA_reg_RNO[63]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[63]_net_1\, D => 
        \sdr_dataout_reg[15]_net_1\, Y => N_201_mux_i);
    
    \sdr_datain_0[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[29]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[13]_net_1\);
    
    \WDATA_reg[55]\ : SLE
      port map(D => \WDATA_mux[55]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[55]_net_1\);
    
    \RDATA_reg_RNO[6]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[6]\, D => 
        \sdr_dataout_reg[6]_net_1\, Y => N_176_mux_i);
    
    \raddr_reg_RNIVU71T[20]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[20]_net_1\, C => 
        \raddr_reg_9_2_axb_20_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_19, S => N_769, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_20);
    
    \RDATA_reg_RNIRICN1[16]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[16]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_2_i_1_0);
    
    \RDATA_reg[56]\ : SLE
      port map(D => N_194_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[56]_net_1\);
    
    \WDATA_mux_3_0[11]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[11]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[11]_net_1\, Y => \WDATA_mux[11]\);
    
    \RDATA_reg_RNITPHN1[63]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[63]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i17_mux_i_1);
    
    \WDATA_reg[12]\ : SLE
      port map(D => \WDATA_mux[12]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[12]_net_1\);
    
    \RDATA_reg_RNO[5]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[5]\, D => 
        \sdr_dataout_reg[5]_net_1\, Y => N_175_mux_i);
    
    \WDATA_mux_3_0_a2_0[7]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \asize_reg[0]_net_1\, B => 
        \asize_reg[1]_net_1\, C => COREAXI_0_AXImslave16_WSTRB(0), 
        D => COREAXI_0_AXImslave16_WSTRB(4), Y => N_3268);
    
    \WDATA_mux_3_0[6]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[6]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[6]_net_1\, Y => \WDATA_mux[6]\);
    
    \RDATA_reg[44]\ : SLE
      port map(D => \sdr_dataout_reg[12]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[44]_net_1\);
    
    \RDATA_reg[15]\ : SLE
      port map(D => N_185_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[15]\);
    
    \WSTRB_reg[3]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(3), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[3]_net_1\);
    
    \sdr_datain_3[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[0]_net_1\, C => \WDATA_reg[0]_net_1\, Y => 
        \sdr_datain_3[0]_net_1\);
    
    \RDATA_reg_RNISOCR1[47]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[15]\, B => 
        \RDATA_reg[47]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_47);
    
    \raddr_reg_9[6]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_755, Y => \raddr_reg_9[6]_net_1\);
    
    \WDATA_reg[40]\ : SLE
      port map(D => \WDATA_mux[40]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[40]_net_1\);
    
    \WDATA_reg_RNO[35]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(35), 
        Y => \WDATA_mux[35]\);
    
    \WDATA_mux_3_0[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(56), B => 
        COREAXI_0_AXImslave16_WDATA(24), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[24]\);
    
    \sdr_count_RNO[1]\ : CFG4
      generic map(INIT => x"006C")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => un1_sdr_count_0_sqmuxa, D => 
        N_3299, Y => N_3279_i);
    
    \WDATA_mux_8_1[6]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[6]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(38), D
         => COREAXI_0_AXImslave16_WDATA(22), Y => 
        \WDATA_mux_8_1[6]_net_1\);
    
    \RDATA_reg[30]\ : SLE
      port map(D => N_3073_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[30]_net_1\);
    
    \axi_state_ns[3]\ : CFG4
      generic map(INIT => x"7530")

      port map(A => N_23, B => N_349, C => \axi_state[1]_net_1\, 
        D => \axi_state_0\, Y => \axi_state_ns[3]_net_1\);
    
    \WDATA_reg[9]\ : SLE
      port map(D => \WDATA_mux[9]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[9]_net_1\);
    
    \axi_state[4]\ : SLE
      port map(D => \axi_state_ns[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_BVALID\);
    
    \sdr_datain_1[10]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[10]_net_1\, C => \WDATA_reg[58]_net_1\, D
         => \WDATA_reg[42]_net_1\, Y => \sdr_datain_1[10]_net_1\);
    
    \DQM_mux_ns[0]\ : CFG4
      generic map(INIT => x"0257")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => N_3154, C
         => N_3145, D => \DQM_mux_ns_1[0]_net_1\, Y => 
        \DQM_mux[0]\);
    
    \RDATA_reg_RNO[9]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[9]\, D => 
        \sdr_dataout_reg[9]_net_1\, Y => N_179_mux_i);
    
    \raddr_reg_9[20]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_769, Y => \raddr_reg_9[20]_net_1\);
    
    \sdr_datain_3[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[6]_net_1\, C => \WDATA_reg[6]_net_1\, Y => 
        \sdr_datain_3[6]_net_1\);
    
    \WDATA_reg_RNO[47]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(47), 
        Y => \WDATA_mux[47]\);
    
    \RDATA_reg_RNI8NFQ1[36]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[4]\, B => 
        \RDATA_reg[36]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3102_i);
    
    \sdr_datain_reg_RNO[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[1]_net_1\, C => \sdr_datain_1[1]_net_1\, Y
         => \sdr_datain[1]\);
    
    \sdr_datain_2[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[4]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[4]_net_1\);
    
    \WDATA_mux_3[20]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(20), C => 
        \WDATA_mux_31[20]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[20]\);
    
    \sdr_datain_reg[7]\ : SLE
      port map(D => \sdr_datain[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(7));
    
    \WSTRB_mux_3_0_a3_1[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \asize_reg[1]_net_1\, B => 
        \asize_reg[0]_net_1\, Y => N_3157);
    
    WDATA_mux_15_m2s2 : CFG2
      generic map(INIT => x"E")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WSTRB(5), Y => WDATA_mux_15_sm0);
    
    \WDATA_reg[47]\ : SLE
      port map(D => \WDATA_mux[47]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[47]_net_1\);
    
    \sdr_datain_1[13]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[13]_net_1\, C => \WDATA_reg[61]_net_1\, D
         => \WDATA_reg[45]_net_1\, Y => \sdr_datain_1[13]_net_1\);
    
    \WDATA_reg[10]\ : SLE
      port map(D => \WDATA_mux[10]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[10]_net_1\);
    
    \RDATA_reg[37]\ : SLE
      port map(D => \sdr_dataout_reg[5]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[37]_net_1\);
    
    \sdr_datain_reg[4]\ : SLE
      port map(D => \sdr_datain[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(4));
    
    \RDATA_reg_RNII6EK1[30]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[30]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_3\, C => N_3141, D => 
        N_3167_i, Y => N_68_mux_i);
    
    \sdr_datain_reg_RNO[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[12]_net_1\, C => \sdr_datain_1[12]_net_1\, 
        Y => \sdr_datain[12]\);
    
    \raddr_reg_RNIC4BFJ[13]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[13]_net_1\, C => 
        \raddr_reg_9_2_axb_13_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_12, S => N_762, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_13);
    
    \WDATA_mux_3_0_a5_1_0[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(6), B => 
        COREAXI_0_AXImslave16_WDATA(48), Y => \WDATA_mux_8_m0[0]\);
    
    \sdr_datain_0[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[21]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[5]_net_1\);
    
    \WDATA_reg[44]\ : SLE
      port map(D => \WDATA_mux[44]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[44]_net_1\);
    
    \WDATA_mux_3_0_RNO[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => COREAXI_0_AXImslave16_WSTRB(0), B => 
        \WDATA_mux_8_3[4]_net_1\, C => \WDATA_mux_8_1[4]_net_1\, 
        Y => \WDATA_mux_8[4]\);
    
    \RDATA_reg_RNO[52]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[52]_net_1\, D => 
        \sdr_dataout_reg[4]_net_1\, Y => N_190_mux_i);
    
    \RDATA_reg[59]\ : SLE
      port map(D => N_197_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[59]_net_1\);
    
    \raddr_reg_RNITI9LB[7]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[7]_net_1\, C => 
        \raddr_reg_9_2_axb_7_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_6, S => N_756, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_7);
    
    \RDATA_reg[34]\ : SLE
      port map(D => \sdr_dataout_reg[2]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[34]_net_1\);
    
    \axi_state_ns[9]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \axi_state[3]_net_1\, B => RW_ACK, C => 
        \axi_state[0]_net_1\, D => N_338, Y => 
        \axi_state_ns[9]_net_1\);
    
    RAS_N : SLE
      port map(D => RAS_N_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RAS_N_c);
    
    \RDATA_reg_RNIN2TQ[57]\ : CFG4
      generic map(INIT => x"7D41")

      port map(A => \RDATA_reg[57]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        m16_1_1_2, Y => i58_mux_0);
    
    \sdr_datain_2[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[0]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_2[0]_net_1\);
    
    raddr_reg_9_2_axb_8_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(9), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(9), Y => 
        \raddr_reg_9_2_axb_8_1\);
    
    \WDATA_reg[23]\ : SLE
      port map(D => \WDATA_mux[23]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[23]_net_1\);
    
    \WDATA_reg[17]\ : SLE
      port map(D => \WDATA_mux[17]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[17]_net_1\);
    
    \axi_count_RNO[0]\ : CFG4
      generic map(INIT => x"0110")

      port map(A => \COREAXI_0_AXImslave16_BVALID\, B => 
        \axi_state[9]_net_1\, C => N_72, D => N_3281, Y => 
        N_3276_i);
    
    \RDATA_reg_RNIK8EK1[31]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[31]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[15]\, C => N_3141, D => 
        N_3167_i, Y => N_67_mux_i);
    
    un7_wstrb_reg_i_a3 : CFG2
      generic map(INIT => x"1")

      port map(A => \WSTRB_reg[2]_net_1\, B => 
        \WSTRB_reg[3]_net_1\, Y => \un7_wstrb_reg_i_a3\);
    
    \RDATA_reg[46]\ : SLE
      port map(D => \sdr_dataout_reg[14]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_reg_3);
    
    \RDATA_reg_RNIOFTB1[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[3]\, Y => N_3170_i);
    
    \WDATA_mux_3_0[9]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_15[9]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[9]_net_1\, Y => \WDATA_mux[9]\);
    
    \RDATA_reg_RNIOGDN1[22]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[22]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_3_i_1_0);
    
    \WDATA_reg_RNO[34]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(34), 
        Y => \WDATA_mux[34]\);
    
    \WDATA_mux_15_3[12]\ : CFG4
      generic map(INIT => x"CACE")

      port map(A => COREAXI_0_AXImslave16_WSTRB(3), B => 
        COREAXI_0_AXImslave16_WDATA(12), C => WDATA_mux_15_sm0, D
         => COREAXI_0_AXImslave16_WSTRB(5), Y => 
        \WDATA_mux_15_3[12]_net_1\);
    
    \sdr_datain_0[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[30]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[14]_net_1\);
    
    \WDATA_mux_3[19]\ : CFG4
      generic map(INIT => x"D844")

      port map(A => \asize_reg[0]_net_1\, B => 
        COREAXI_0_AXImslave16_WDATA(19), C => 
        \WDATA_mux_31[19]_net_1\, D => \asize_reg[1]_net_1\, Y
         => \WDATA_mux[19]\);
    
    \un1_B_SIZE_reg_0_a2[2]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \B_SIZE_reg[0]_net_1\, B => N_335_i, C => 
        N_343_i, Y => \un1_B_SIZE_reg_0_a2[2]_net_1\);
    
    \WDATA_mux_3_0_RNO[9]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \WDATA_mux_15_3[9]_net_1\, B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        \WDATA_mux_15_1[9]_net_1\, Y => \WDATA_mux_15[9]\);
    
    \RDATA_reg_RNINFDN1[21]\ : CFG4
      generic map(INIT => x"3313")

      port map(A => \RDATA_reg[21]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_4_i_1_0);
    
    \WDATA_reg[14]\ : SLE
      port map(D => \WDATA_mux[14]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[14]_net_1\);
    
    \WDATA_mux_15_1[11]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[11]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(27), D
         => COREAXI_0_AXImslave16_WDATA(43), Y => 
        \WDATA_mux_15_1[11]_net_1\);
    
    \RDATA_reg[6]\ : SLE
      port map(D => N_176_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA[6]\);
    
    \WDATA_mux_8_0[0]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8_m0[0]\, B => 
        COREAXI_0_AXImslave16_WSTRB(4), C => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_8_0[0]_net_1\);
    
    \RDATA_reg_RNO[1]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[1]\, D => 
        \sdr_dataout_reg[1]_net_1\, Y => N_171_mux_i);
    
    \RDATA_reg_RNO[0]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[0]\, D => 
        \sdr_dataout_reg[0]_net_1\, Y => N_170_mux_i);
    
    asize_reg_134 : CFG3
      generic map(INIT => x"CA")

      port map(A => \asize_reg[0]_net_1\, B => \asize[0]_net_1\, 
        C => N_295_i, Y => \asize_reg_134\);
    
    \WSTRB_reg[1]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(1), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[1]_net_1\);
    
    \WDATA_reg[7]\ : SLE
      port map(D => \WDATA_mux[7]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[7]_net_1\);
    
    \raddr_reg_9[10]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_759, Y => \raddr_reg_9[10]_net_1\);
    
    \sdr_datain_reg_RNO[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[4]_net_1\, C => \sdr_datain_1[4]_net_1\, Y
         => \sdr_datain[4]\);
    
    raddr_reg_9_2_axb_3_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(4), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(4), Y => 
        \raddr_reg_9_2_axb_3_1\);
    
    \RDATA_reg_RNO[13]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => 
        \COREAXI_0_AXImslave16_RDATA[13]\, D => 
        \sdr_dataout_reg[13]_net_1\, Y => N_183_mux_i);
    
    \RDATA_reg[21]\ : SLE
      port map(D => \sdr_dataout_reg[5]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[19]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[21]_net_1\);
    
    \sdr_datain_3[5]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[5]_net_1\, C => \WDATA_reg[5]_net_1\, Y => 
        \sdr_datain_3[5]_net_1\);
    
    \axi_state_ns_0_o2[7]\ : CFG3
      generic map(INIT => x"FD")

      port map(A => \axi_count[0]_net_1\, B => N_3286, C => 
        \axi_count[3]_net_1\, Y => \N_3297\);
    
    \RDATA_reg_RNI6DHJ1[23]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[23]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[7]\, C => N_3141, D => 
        N_3167_i, Y => COREAXI_0_AXImslave16_RDATA_m_23);
    
    \raddr_reg_RNIEOL0E[9]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[9]_net_1\, C => 
        \raddr_reg_9_2_axb_9_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_8, S => N_758, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_9);
    
    \WDATA_mux_3_0[31]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(63), B => 
        COREAXI_0_AXImslave16_WDATA(31), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[31]\);
    
    \RDATA_reg[55]\ : SLE
      port map(D => N_193_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[55]_net_1\);
    
    CAS_N : SLE
      port map(D => CAS_N_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => CAS_N_c);
    
    \WSTRB_reg[0]\ : SLE
      port map(D => COREAXI_0_AXImslave16_WSTRB(0), CLK => 
        SDRCLK_c, EN => \WREADY_SI16\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WSTRB_reg[0]_net_1\);
    
    \sdr_datain_0[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \WDATA_reg[20]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \sdr_count[1]_net_1\, Y => 
        \sdr_datain_0[4]_net_1\);
    
    \WDATA_mux_3_0_a5_2[14]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => COREAXI_0_AXImslave16_WDATA(46), B => 
        COREAXI_0_AXImslave16_WSTRB(1), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => N_3157, Y => N_3202);
    
    \RDATA_reg_RNI2HFQ1[33]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[1]\, B => 
        \RDATA_reg[33]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_33);
    
    \xhdl21.b_size4\ : CFG2
      generic map(INIT => x"4")

      port map(A => \asize[1]_net_1\, B => \asize[0]_net_1\, Y
         => b_size4);
    
    \WDATA_mux_8_3[0]\ : CFG4
      generic map(INIT => x"E2F2")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(0), D
         => COREAXI_0_AXImslave16_WSTRB(4), Y => 
        \WDATA_mux_8_3[0]_net_1\);
    
    \WDATA_reg[32]\ : SLE
      port map(D => \WDATA_mux[32]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[32]_net_1\);
    
    \WDATA_mux_15_0[8]\ : CFG4
      generic map(INIT => x"FF08")

      port map(A => COREAXI_0_AXImslave16_WDATA(56), B => 
        COREAXI_0_AXImslave16_WSTRB(7), C => 
        COREAXI_0_AXImslave16_WSTRB(5), D => 
        COREAXI_0_AXImslave16_WSTRB(3), Y => 
        \WDATA_mux_15_0[8]_net_1\);
    
    \WSTRB_mux_3_0_a3[0]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \WSTRB_reg[1]_net_1\, B => 
        \WSTRB_reg[4]_net_1\, C => \un7_wstrb_reg_i_a3\, D => 
        N_3157, Y => N_3154);
    
    \WDATA_reg_RNO[53]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(53), 
        Y => \WDATA_mux[53]\);
    
    \RDATA_reg_RNO[30]\ : CFG4
      generic map(INIT => x"F2D0")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[30]_net_1\, D => 
        \sdr_dataout_reg[14]_net_1\, Y => N_3073_i);
    
    \RDATA_reg_RNO[61]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[61]_net_1\, D => 
        \sdr_dataout_reg[13]_net_1\, Y => N_199_mux_i);
    
    raddr_reg_9_2_axb_21_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(22), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(22), Y => 
        \raddr_reg_9_2_axb_21_1\);
    
    \RDATA_reg_RNI8FHJ1[24]\ : CFG4
      generic map(INIT => x"00AC")

      port map(A => \RDATA_reg[24]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA[8]\, C => N_3141, D => 
        N_3167_i, Y => N_79_mux_i);
    
    \RDATA_reg_RNIMDTB1[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[1]\, Y => 
        COREAXI_0_AXImslave16_RDATA_m_1);
    
    \WDATA_reg[46]\ : SLE
      port map(D => \WDATA_mux[46]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[46]_net_1\);
    
    \SA[5]\ : SLE
      port map(D => \SA_i[5]\, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => SA_c(5));
    
    \sdr_datain_3[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_2[3]_net_1\, C => \WDATA_reg[3]_net_1\, Y => 
        \sdr_datain_3[3]_net_1\);
    
    \sdr_datain_reg_RNO[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[8]_net_1\, C => \sdr_datain_1[8]_net_1\, Y
         => \sdr_datain[8]\);
    
    \sdr_datain_1[14]\ : CFG4
      generic map(INIT => x"E6C4")

      port map(A => \sdr_count[1]_net_1\, B => 
        \sdr_datain_0[14]_net_1\, C => \WDATA_reg[62]_net_1\, D
         => \WDATA_reg[46]_net_1\, Y => \sdr_datain_1[14]_net_1\);
    
    \RDATA_reg_RNIQ4HH[19]\ : CFG4
      generic map(INIT => x"0530")

      port map(A => \COREAXI_0_AXImslave16_RDATA[3]\, B => 
        \RDATA_reg[19]_net_1\, C => \asize_reg[1]_net_1\, D => 
        \asize_reg[0]_net_1\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_i_0[51]\);
    
    \RDATA_regce[19]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \sdr_count[1]_net_1\, B => \R_VALID\, C => 
        \sdr_count[0]_net_1\, Y => \RDATA_regce[19]_net_1\);
    
    \RDATA_reg[36]\ : SLE
      port map(D => \sdr_dataout_reg[4]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[36]_net_1\);
    
    \sdr_dataout_reg[14]\ : SLE
      port map(D => DQ_in(14), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[14]_net_1\);
    
    \sdr_datain_reg_RNO[9]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \sdr_count_RNI201B[3]_net_1\, B => 
        \sdr_datain_3[9]_net_1\, C => \sdr_datain_1[9]_net_1\, Y
         => \sdr_datain[9]\);
    
    \WDATA_reg[51]\ : SLE
      port map(D => \WDATA_mux[51]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[51]_net_1\);
    
    \RDATA_reg[49]\ : SLE
      port map(D => N_187_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_reg[49]_net_1\);
    
    axi_nextstate_1_sqmuxa_i_o2_i_a2_i : CFG3
      generic map(INIT => x"BF")

      port map(A => \N_389\, B => COREAXI_0_AXImslave16_WVALID, C
         => \axi_state[5]_net_1\, Y => WREADY_SI16_i);
    
    \RDATA_reg_RNISJTB1[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_3167_i, B => 
        \COREAXI_0_AXImslave16_RDATA[7]\, Y => 
        \COREAXI_0_AXImslave16_RDATA_m_7\);
    
    \raddr_reg_9[9]\ : CFG4
      generic map(INIT => x"FB00")

      port map(A => COREAXI_0_AXImslave16_AWVALID, B => 
        \axi_state[9]_net_1\, C => COREAXI_0_AXImslave16_ARVALID, 
        D => N_758, Y => \raddr_reg_9[9]_net_1\);
    
    \WDATA_reg[5]\ : SLE
      port map(D => \WDATA_mux[5]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[5]_net_1\);
    
    \sdr_datain_reg[14]\ : SLE
      port map(D => \sdr_datain[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sdr_datain_reg(14));
    
    \WDATA_mux_15_1[10]\ : CFG4
      generic map(INIT => x"E6A2")

      port map(A => \WDATA_mux_15_0[10]_net_1\, B => 
        WDATA_mux_15_sm0, C => COREAXI_0_AXImslave16_WDATA(26), D
         => COREAXI_0_AXImslave16_WDATA(42), Y => 
        \WDATA_mux_15_1[10]_net_1\);
    
    \WDATA_reg[61]\ : SLE
      port map(D => \WDATA_mux[61]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[61]_net_1\);
    
    \RDATA_reg_RNO[58]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[58]_net_1\, D => 
        \sdr_dataout_reg[10]_net_1\, Y => N_196_mux_i);
    
    \RDATA_reg_RNIQMHN1[60]\ : CFG4
      generic map(INIT => x"3CBE")

      port map(A => \RDATA_reg[60]_net_1\, B => 
        \asize_reg[0]_net_1\, C => \asize_reg[1]_net_1\, D => 
        N_3167_i, Y => i22_mux_i_1);
    
    \RDATA_reg[11]\ : SLE
      port map(D => N_181_mux_i, CLK => SDRCLK_c, EN => \R_VALID\, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAXI_0_AXImslave16_RDATA_0\);
    
    \WDATA_mux_31[17]\ : CFG4
      generic map(INIT => x"CCA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(49), B => 
        COREAXI_0_AXImslave16_WDATA(17), C => 
        COREAXI_0_AXImslave16_WSTRB(6), D => 
        COREAXI_0_AXImslave16_WSTRB(2), Y => 
        \WDATA_mux_31[17]_net_1\);
    
    \asize_reg_RNI28505[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_4\, C => i22_mux_5_i_1_0, 
        D => i22_mux_5_i_1, Y => i22_mux_5_i);
    
    \WDATA_reg[16]\ : SLE
      port map(D => \WDATA_mux[16]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[16]_net_1\);
    
    \WDATA_reg_RNO[59]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(59), 
        Y => \WDATA_mux[59]\);
    
    \WDATA_reg[30]\ : SLE
      port map(D => \WDATA_mux[30]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[30]_net_1\);
    
    \asize_reg_RNIBH505[1]\ : CFG4
      generic map(INIT => x"5E00")

      port map(A => \asize_reg[1]_net_1\, B => 
        \COREAXI_0_AXImslave16_RDATA_m_7\, C => i22_mux_2_i_1_0, 
        D => i22_mux_2_i_1, Y => i22_mux_2_i);
    
    \WDATA_reg_RNO[42]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \N_74\, B => COREAXI_0_AXImslave16_WDATA(42), 
        Y => \WDATA_mux[42]\);
    
    \WSTRB_mux_3_0_a3_0_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \WSTRB_reg[3]_net_1\, B => 
        \WSTRB_reg[6]_net_1\, Y => 
        \WSTRB_mux_3_0_a3_0_0[2]_net_1\);
    
    \RDATA_reg_RNIVAN32[49]\ : CFG2
      generic map(INIT => x"1")

      port map(A => N_3167_i, B => i58_mux_2, Y => 
        COREAXI_0_AXImslave16_RDATA_m_49);
    
    \sdr_count[3]\ : SLE
      port map(D => N_3277_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_count[3]_net_1\);
    
    \raddr_reg_9_RNO_0[22]\ : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(23), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(23), Y => 
        raddr_reg_9_2_axb_22_1);
    
    \WDATA_mux_3_0_0[15]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => COREAXI_0_AXImslave16_WDATA(15), B => 
        COREAXI_0_AXImslave16_WDATA(47), C => N_3210, D => N_3236, 
        Y => \WDATA_mux_3_0_0[15]_net_1\);
    
    \sdr_dataout_reg[9]\ : SLE
      port map(D => DQ_in(9), CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sdr_dataout_reg[9]_net_1\);
    
    \RDATA_reg_RNO[50]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => \sdr_count[0]_net_1\, B => 
        \sdr_count[1]_net_1\, C => \RDATA_reg[50]_net_1\, D => 
        \sdr_dataout_reg[2]_net_1\, Y => N_188_mux_i);
    
    \RDATA_reg_RNIKQ192[51]\ : CFG4
      generic map(INIT => x"0504")

      port map(A => \COREAXI_0_AXImslave16_RDATA_m_i_0[51]\, B
         => \RDATA_reg[51]_net_1\, C => N_3167_i, D => \N_74\, Y
         => N_8_i);
    
    asize_reg_135 : CFG3
      generic map(INIT => x"3A")

      port map(A => \asize_reg[1]_net_1\, B => \asize[1]_net_1\, 
        C => N_295_i, Y => \asize_reg_135\);
    
    \DQM_mux_ns_1_1[1]\ : CFG3
      generic map(INIT => x"1D")

      port map(A => \WSTRB_reg[5]_net_1\, B => 
        \sdr_count[0]_net_1\, C => \WSTRB_reg[7]_net_1\, Y => 
        \DQM_mux_ns_1_1[1]_net_1\);
    
    \un7_1.SUM_i_o2[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => N_3281, B => \axi_count[0]_net_1\, Y => 
        N_3289);
    
    \WDATA_reg[37]\ : SLE
      port map(D => \WDATA_mux[37]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[37]_net_1\);
    
    \WDATA_mux_3_0[2]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[2]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[2]_net_1\, Y => \WDATA_mux[2]\);
    
    \RDATA_reg[45]\ : SLE
      port map(D => \sdr_dataout_reg[13]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[45]_net_1\);
    
    \raddr_reg_RNI3N0RK[14]\ : ARI1
      generic map(INIT => x"4A300")

      port map(A => VCC_net_1, B => \raddr_reg[14]_net_1\, C => 
        \raddr_reg_9_2_axb_14_1\, D => raddr_reg_9_sn_N_3_i, FCI
         => raddr_reg_9_2_cry_13, S => N_763, Y => OPEN, FCO => 
        raddr_reg_9_2_cry_14);
    
    \RDATA_reg_RNIAPFQ1[37]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \COREAXI_0_AXImslave16_RDATA[5]\, B => 
        \RDATA_reg[37]_net_1\, C => N_3167_i, D => \N_74\, Y => 
        N_3100_i);
    
    \WDATA_reg[49]\ : SLE
      port map(D => \WDATA_mux[49]\, CLK => SDRCLK_c, EN => 
        \WREADY_SI16\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_reg[49]_net_1\);
    
    \WDATA_mux_8_1[4]\ : CFG4
      generic map(INIT => x"EA62")

      port map(A => \WDATA_mux_8_0[4]_net_1\, B => 
        WDATA_mux_8_sm0, C => COREAXI_0_AXImslave16_WDATA(36), D
         => COREAXI_0_AXImslave16_WDATA(20), Y => 
        \WDATA_mux_8_1[4]_net_1\);
    
    \WDATA_mux_3_0[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => COREAXI_0_AXImslave16_WDATA(61), B => 
        COREAXI_0_AXImslave16_WDATA(29), C => N_3172, D => N_3207, 
        Y => \WDATA_mux[29]\);
    
    raddr_reg_9_2_axb_6_1 : CFG3
      generic map(INIT => x"47")

      port map(A => COREAXI_0_AXImslave16_ARADDR(7), B => 
        COREAXI_0_AXImslave16_ARVALID, C => 
        COREAXI_0_AXImslave16_AWADDR(7), Y => 
        \raddr_reg_9_2_axb_6_1\);
    
    \RDATA_reg[39]\ : SLE
      port map(D => \sdr_dataout_reg[7]_net_1\, CLK => SDRCLK_c, 
        EN => \RDATA_regce[32]_net_1\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RDATA_reg[39]_net_1\);
    
    WDATA_mux_8_m2s2 : CFG2
      generic map(INIT => x"E")

      port map(A => COREAXI_0_AXImslave16_WSTRB(2), B => 
        COREAXI_0_AXImslave16_WSTRB(4), Y => WDATA_mux_8_sm0);
    
    \WDATA_mux_3_0[0]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \WDATA_mux_8[0]\, B => N_3141, C => 
        \WDATA_mux_3_0_0[0]_net_1\, Y => \WDATA_mux[0]\);
    
    \raddr_reg[3]\ : SLE
      port map(D => \raddr_reg_9[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_reg[3]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( top_sb_0_POWER_ON_RESET_N             : in    std_logic;
          top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic;
          top_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic;
          CORERESETP_0_RESET_N_F2M              : out   std_logic;
          SDRCLK_c                              : in    std_logic;
          MSS_READY                             : out   std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \MSS_HPMS_READY_int\, \mss_ready_select\, VCC_net_1, 
        \sm1_areset_n_clk_base\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, GND_net_1, 
        \mss_ready_state\, \RESET_N_M2F_clk_base\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_clk_base\, 
        \FIC_2_APB_M_PRESET_N_q1\, sm1_areset_n_q1, 
        \MSS_HPMS_READY_int_3\ : std_logic;

begin 


    MSS_HPMS_READY_int_RNI5MMF : CLKINT
      port map(A => \MSS_HPMS_READY_int\, Y => MSS_READY);
    
    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => top_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RESET_N_M2F_clk_base\);
    
    RESET_N_F2M_int : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => \sm1_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORERESETP_0_RESET_N_F2M);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => 
        \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \sm1_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    sm1_areset_n_clk_base : SLE
      port map(D => sm1_areset_n_q1, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => top_sb_0_POWER_ON_RESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm1_areset_n_clk_base\);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => 
        \RESET_N_M2F_clk_base\, ALn => \sm1_areset_n_clk_base\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mss_ready_state\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => top_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_q1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \FIC_2_APB_M_PRESET_N_clk_base\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => top_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        sm1_areset_n_q1);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => \sm1_areset_n_clk_base\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \MSS_HPMS_READY_int\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVEARBITER_1 is

    port( masterAddrInProg                           : out   std_logic_vector(3 downto 0);
          current_state_0                            : in    std_logic;
          xhdl1221_0                                 : in    std_logic;
          regHMASTLOCK                               : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK : in    std_logic;
          masterRegAddrSel                           : in    std_logic;
          SDRCLK_c                                   : in    std_logic;
          MSS_READY                                  : in    std_logic
        );

end COREAHBLITE_SLAVEARBITER_1;

architecture DEF_ARCH of COREAHBLITE_SLAVEARBITER_1 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \arbRegSMCurrentState[1]_net_1\, VCC_net_1, N_141_i, 
        GND_net_1, \masterAddrInProg[3]\, N_143_i, 
        \arbRegSMCurrentState[15]_net_1\, N_119_i, 
        \arbRegSMCurrentState[14]_net_1\, N_121_i, 
        \arbRegSMCurrentState[13]_net_1\, N_123_i, 
        \arbRegSMCurrentState[12]_net_1\, N_125_i, 
        \arbRegSMCurrentState[10]_net_1\, 
        \arbRegSMCurrentState_ns[5]_net_1\, 
        \arbRegSMCurrentState[9]_net_1\, N_129_i, 
        \masterAddrInProg[1]\, N_131_i, 
        \arbRegSMCurrentState[6]_net_1\, 
        \arbRegSMCurrentState_ns[9]_net_1\, 
        \arbRegSMCurrentState[5]_net_1\, N_135_i, 
        \masterAddrInProg[2]\, N_137_i, 
        \arbRegSMCurrentState[2]_net_1\, 
        \arbRegSMCurrentState_ns[13]_net_1\, N_4_0, N_148_0, 
        N_5_0, N_69, N_148, \arbRegSMCurrentState_ns_i_0_a2_0[1]\, 
        N_94, N_170, N_146, 
        \arbRegSMCurrentState_ns_i_0_a2_1_0[2]_net_1\, N_101, 
        N_68, \arbRegSMCurrentState_ns_i_0_0[1]_net_1\, 
        \arbRegSMCurrentState_ns_i_0_1[2]_net_1\ : std_logic;

begin 

    masterAddrInProg(3) <= \masterAddrInProg[3]\;
    masterAddrInProg(2) <= \masterAddrInProg[2]\;
    masterAddrInProg(1) <= \masterAddrInProg[1]\;

    \arbRegSMCurrentState_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => current_state_0, B => \masterAddrInProg[3]\, 
        Y => N_141_i);
    
    \arbRegSMCurrentState_ns_i_0_a2_3[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \arbRegSMCurrentState[2]_net_1\, B => 
        \arbRegSMCurrentState[14]_net_1\, C => 
        \arbRegSMCurrentState[10]_net_1\, D => 
        \arbRegSMCurrentState[6]_net_1\, Y => N_148);
    
    \arbRegSMCurrentState_RNIUIKV[13]\ : CFG3
      generic map(INIT => x"2E")

      port map(A => N_148_0, B => N_4_0, C => 
        \arbRegSMCurrentState[13]_net_1\, Y => N_5_0);
    
    \arbRegSMCurrentState_ns[13]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[1]_net_1\, B => 
        \arbRegSMCurrentState[2]_net_1\, C => xhdl1221_0, Y => 
        \arbRegSMCurrentState_ns[13]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_a2_1[1]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \arbRegSMCurrentState[13]_net_1\, B => 
        xhdl1221_0, C => \arbRegSMCurrentState[14]_net_1\, D => 
        \arbRegSMCurrentState[15]_net_1\, Y => N_101);
    
    \arbRegSMCurrentState[12]\ : SLE
      port map(D => N_125_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[12]_net_1\);
    
    \arbRegSMCurrentState_ns[9]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[5]_net_1\, B => 
        \arbRegSMCurrentState[6]_net_1\, C => xhdl1221_0, Y => 
        \arbRegSMCurrentState_ns[9]_net_1\);
    
    \arbRegSMCurrentState[8]\ : SLE
      port map(D => N_131_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[1]\);
    
    \arbRegSMCurrentState[10]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[5]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \arbRegSMCurrentState[10]_net_1\);
    
    g0_3_m4_0 : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, C => 
        regHMASTLOCK, Y => N_4_0);
    
    \arbRegSMCurrentState_RNI6QK5[2]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \arbRegSMCurrentState[2]_net_1\, B => 
        \arbRegSMCurrentState[14]_net_1\, C => 
        \arbRegSMCurrentState[10]_net_1\, D => 
        \arbRegSMCurrentState[6]_net_1\, Y => N_148_0);
    
    \arbRegSMCurrentState_ns_i_0_a2_2[2]\ : CFG4
      generic map(INIT => x"010B")

      port map(A => masterRegAddrSel, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, C => 
        \arbRegSMCurrentState[12]_net_1\, D => regHMASTLOCK, Y
         => N_170);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \arbRegSMCurrentState_RNO[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => current_state_0, B => \masterAddrInProg[3]\, 
        Y => N_143_i);
    
    \arbRegSMCurrentState[0]\ : SLE
      port map(D => N_143_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[3]\);
    
    \arbRegSMCurrentState_RNO[12]\ : CFG4
      generic map(INIT => x"0A0E")

      port map(A => \arbRegSMCurrentState[12]_net_1\, B => 
        \arbRegSMCurrentState[13]_net_1\, C => current_state_0, D
         => N_94, Y => N_125_i);
    
    \arbRegSMCurrentState_RNO[15]\ : CFG4
      generic map(INIT => x"0045")

      port map(A => current_state_0, B => 
        \arbRegSMCurrentState[15]_net_1\, C => N_68, D => N_146, 
        Y => N_119_i);
    
    \arbRegSMCurrentState_RNO[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => current_state_0, B => \masterAddrInProg[1]\, 
        Y => N_131_i);
    
    \arbRegSMCurrentState[14]\ : SLE
      port map(D => N_121_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[14]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_o2[3]\ : CFG4
      generic map(INIT => x"47FF")

      port map(A => regHMASTLOCK, B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, D => 
        xhdl1221_0, Y => N_94);
    
    \arbRegSMCurrentState[6]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[9]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \arbRegSMCurrentState[6]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_o2[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => xhdl1221_0, B => 
        \arbRegSMCurrentState[14]_net_1\, Y => N_69);
    
    \arbRegSMCurrentState[1]\ : SLE
      port map(D => N_141_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \arbRegSMCurrentState_RNIBMJN3[12]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => N_5_0, B => xhdl1221_0, C => 
        \arbRegSMCurrentState[12]_net_1\, D => 
        \arbRegSMCurrentState[15]_net_1\, Y => 
        masterAddrInProg(0));
    
    \arbRegSMCurrentState_RNO[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => current_state_0, B => \masterAddrInProg[2]\, 
        Y => N_137_i);
    
    \arbRegSMCurrentState_ns_i_0_a2_0[0]\ : CFG4
      generic map(INIT => x"0E04")

      port map(A => masterRegAddrSel, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, C => 
        \arbRegSMCurrentState[15]_net_1\, D => regHMASTLOCK, Y
         => N_146);
    
    \arbRegSMCurrentState_RNO[13]\ : CFG4
      generic map(INIT => x"0E0F")

      port map(A => \arbRegSMCurrentState[13]_net_1\, B => 
        \arbRegSMCurrentState[12]_net_1\, C => 
        \arbRegSMCurrentState_ns_i_0_1[2]_net_1\, D => N_68, Y
         => N_123_i);
    
    \arbRegSMCurrentState_ns_i_0_1[2]\ : CFG4
      generic map(INIT => x"FFAC")

      port map(A => \arbRegSMCurrentState_ns_i_0_a2_1_0[2]_net_1\, 
        B => \arbRegSMCurrentState_ns_i_0_a2_0[1]\, C => 
        xhdl1221_0, D => N_170, Y => 
        \arbRegSMCurrentState_ns_i_0_1[2]_net_1\);
    
    \arbRegSMCurrentState_RNO[14]\ : CFG4
      generic map(INIT => x"010F")

      port map(A => N_146, B => 
        \arbRegSMCurrentState_ns_i_0_a2_0[1]\, C => 
        \arbRegSMCurrentState_ns_i_0_0[1]_net_1\, D => N_69, Y
         => N_121_i);
    
    \arbRegSMCurrentState[9]\ : SLE
      port map(D => N_129_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[9]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_a2_1_0[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_148, B => current_state_0, Y => 
        \arbRegSMCurrentState_ns_i_0_a2_1_0[2]_net_1\);
    
    \arbRegSMCurrentState[4]\ : SLE
      port map(D => N_137_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \masterAddrInProg[2]\);
    
    \arbRegSMCurrentState[13]\ : SLE
      port map(D => N_123_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[13]_net_1\);
    
    \arbRegSMCurrentState[2]\ : SLE
      port map(D => \arbRegSMCurrentState_ns[13]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \arbRegSMCurrentState[2]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_o2[2]\ : CFG2
      generic map(INIT => x"D")

      port map(A => xhdl1221_0, B => N_148, Y => N_68);
    
    \arbRegSMCurrentState[5]\ : SLE
      port map(D => N_135_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[5]_net_1\);
    
    \arbRegSMCurrentState_ns_i_0_0[1]\ : CFG4
      generic map(INIT => x"FF10")

      port map(A => \arbRegSMCurrentState[15]_net_1\, B => 
        \arbRegSMCurrentState[13]_net_1\, C => N_148, D => N_101, 
        Y => \arbRegSMCurrentState_ns_i_0_0[1]_net_1\);
    
    \arbRegSMCurrentState[15]\ : SLE
      port map(D => N_119_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \arbRegSMCurrentState[15]_net_1\);
    
    \arbRegSMCurrentState_ns[5]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \arbRegSMCurrentState[9]_net_1\, B => 
        \arbRegSMCurrentState[10]_net_1\, C => xhdl1221_0, Y => 
        \arbRegSMCurrentState_ns[5]_net_1\);
    
    \arbRegSMCurrentState_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => current_state_0, B => \masterAddrInProg[2]\, 
        Y => N_135_i);
    
    \arbRegSMCurrentState_RNO[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => current_state_0, B => \masterAddrInProg[1]\, 
        Y => N_129_i);
    
    \arbRegSMCurrentState_ns_i_0_a2_0_0[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => current_state_0, B => 
        \arbRegSMCurrentState[13]_net_1\, Y => 
        \arbRegSMCurrentState_ns_i_0_a2_0[1]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_SLAVESTAGE_0 is

    port( CoreAHBLite_0_AHBmslave10_HADDR             : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 0);
          regHADDR                                    : in    std_logic_vector(27 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE             : out   std_logic_vector(1 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE  : in    std_logic_vector(1 downto 0);
          regHSIZE                                    : in    std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA            : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0);
          xhdl1221_0                                  : in    std_logic;
          masterAddrInProg_0                          : out   std_logic;
          xhdl1292_0                                  : out   std_logic;
          xhdl1222_0                                  : in    std_logic;
          current_state_0                             : in    std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK         : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK  : in    std_logic;
          masterRegAddrSel                            : in    std_logic;
          regHMASTLOCK                                : in    std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE            : out   std_logic;
          N_91                                        : in    std_logic;
          hsel2                                       : out   std_logic;
          hsel2_0_a2_1                                : out   std_logic;
          SDRCLK_c                                    : in    std_logic;
          MSS_READY                                   : in    std_logic
        );

end COREAHBLITE_SLAVESTAGE_0;

architecture DEF_ARCH of COREAHBLITE_SLAVESTAGE_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVEARBITER_1
    port( masterAddrInProg                           : out   std_logic_vector(3 downto 0);
          current_state_0                            : in    std_logic := 'U';
          xhdl1221_0                                 : in    std_logic := 'U';
          regHMASTLOCK                               : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK : in    std_logic := 'U';
          masterRegAddrSel                           : in    std_logic := 'U';
          SDRCLK_c                                   : in    std_logic := 'U';
          MSS_READY                                  : in    std_logic := 'U'
        );
  end component;

    signal \masterDataInProg[0]_net_1\, VCC_net_1, 
        \masterDataInProg_90\, GND_net_1, 
        \masterDataInProg[1]_net_1\, \masterAddrInProg[1]\, 
        \masterDataInProg[2]_net_1\, \masterAddrInProg[2]\, 
        \masterDataInProg[3]_net_1\, \masterAddrInProg[3]\, 
        hsel2_0_a2_1_net_1, \hwdata10\, \masterAddrInProg_0\, 
        \hsel2\ : std_logic;

    for all : COREAHBLITE_SLAVEARBITER_1
	Use entity work.COREAHBLITE_SLAVEARBITER_1(DEF_ARCH);
begin 

    masterAddrInProg_0 <= \masterAddrInProg_0\;
    hsel2 <= \hsel2\;
    hsel2_0_a2_1 <= hsel2_0_a2_1_net_1;

    \masterDataInProg[3]\ : SLE
      port map(D => \masterAddrInProg[3]\, CLK => SDRCLK_c, EN
         => current_state_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \masterDataInProg[3]_net_1\);
    
    hwdata10_RNILBHG_29 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(1));
    
    \hsel2_0_a2_1\ : CFG3
      generic map(INIT => x"01")

      port map(A => \masterAddrInProg[3]\, B => 
        \masterAddrInProg[2]\, C => \masterAddrInProg[1]\, Y => 
        hsel2_0_a2_1_net_1);
    
    hwdata10_RNILBHG_24 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(6));
    
    hwdata10_RNILBHG_23 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(7));
    
    hsel2_0_a2_RNIQUVN : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(2), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(2));
    
    hwdata10_RNILBHG_28 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(2));
    
    hwdata10_RNILBHG_11 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(19));
    
    hsel2_0_a2_RNIRVVN : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(3), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(3));
    
    hwdata10_RNILBHG_26 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(4));
    
    hsel2_0_a2_RNIAK2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(20), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(20));
    
    hwdata10_RNILBHG_1 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(29));
    
    hsel2_0_a2_RNIPK2Q : CFG4
      generic map(INIT => x"B800")

      port map(A => regHSIZE(1), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HSIZE(1));
    
    hsel2_0_a2_RNIEO2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(24), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(24));
    
    hwdata10_RNILBHG_9 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(21));
    
    hsel2_0_a2_RNIHR2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(27), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(27));
    
    hwdata10_RNILBHG_20 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(10));
    
    hsel2_0_a2_RNIJA9V : CFG4
      generic map(INIT => x"B800")

      port map(A => regHMASTLOCK, B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, D => \hsel2\, 
        Y => CoreAHBLite_0_AHBmslave10_HMASTLOCK);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    hwdata10_RNILBHG_22 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(8));
    
    hsel2_0_a2_RNIFP2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(25), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(25));
    
    hsel2_0_a2_RNI9I1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(10), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(10));
    
    hsel2_0_a2_RNIGP1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(17), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(17));
    
    hwdata10_RNILBHG_25 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(5));
    
    \masterDataInProg[2]\ : SLE
      port map(D => \masterAddrInProg[2]\, CLK => SDRCLK_c, EN
         => current_state_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \masterDataInProg[2]_net_1\);
    
    hwdata10_RNILBHG_0 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(30));
    
    hwdata10_RNILBHG : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(31));
    
    hsel2_0_a2_RNIDN2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(23), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(23));
    
    hsel2_0_a2_RNIOSVN : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(0), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(0));
    
    hsel2_0_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => \masterAddrInProg_0\, B => hsel2_0_a2_1_net_1, 
        Y => \hsel2\);
    
    hsel2_0_a2_RNIPTVN : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(1), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(1));
    
    hsel2_0_a2_1_RNI4J454 : CFG3
      generic map(INIT => x"80")

      port map(A => \masterAddrInProg_0\, B => hsel2_0_a2_1_net_1, 
        C => N_91, Y => CoreAHBLite_0_AHBmslave10_HWRITE);
    
    hwdata10_RNILBHG_17 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(13));
    
    hsel2_0_a2_RNIFO1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(16), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(16));
    
    hwdata10_RNILBHG_5 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(25));
    
    hwdata10_RNILBHG_19 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(11));
    
    hsel2_0_a2_RNIOJ2Q : CFG4
      generic map(INIT => x"B800")

      port map(A => regHSIZE(0), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HSIZE(0));
    
    hwdata10_RNILBHG_3 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(27));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    hsel2_0_a2_RNIV30O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(7), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(7));
    
    \masterDataInProg[1]\ : SLE
      port map(D => \masterAddrInProg[1]\, CLK => SDRCLK_c, EN
         => current_state_0, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \masterDataInProg[1]_net_1\);
    
    \masterDataInProg[0]\ : SLE
      port map(D => \masterDataInProg_90\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \masterDataInProg[0]_net_1\);
    
    hwdata10_RNILBHG_6 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(24));
    
    hsel2_0_a2_RNI050O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(8), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(8));
    
    \MDATAREADY_5_iv[0]\ : CFG3
      generic map(INIT => x"D5")

      port map(A => xhdl1222_0, B => current_state_0, C => 
        \masterDataInProg[0]_net_1\, Y => xhdl1292_0);
    
    hwdata10_RNILBHG_14 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(16));
    
    hwdata10_RNILBHG_13 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(17));
    
    masterDataInProg_90 : CFG3
      generic map(INIT => x"D8")

      port map(A => current_state_0, B => \masterAddrInProg_0\, C
         => \masterDataInProg[0]_net_1\, Y => 
        \masterDataInProg_90\);
    
    hwdata10_RNILBHG_18 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(12));
    
    hsel2_0_a2_RNIIR1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(19), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(19));
    
    hwdata10_RNILBHG_16 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(14));
    
    hsel2_0_a2_RNIBL2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(21), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(21));
    
    hwdata10_RNILBHG_4 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(26));
    
    hsel2_0_a2_RNI160O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(9), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(9));
    
    hsel2_0_a2_RNIDM1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(14), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(14));
    
    hwdata10_RNILBHG_10 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(20));
    
    hwdata10_RNILBHG_21 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(9));
    
    hwdata10_RNILBHG_12 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(18));
    
    hsel2_0_a2_RNICM2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(22), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(22));
    
    hwdata10_RNILBHG_15 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(15));
    
    hwdata10_RNILBHG_2 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(28));
    
    hsel2_0_a2_RNIHQ1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(18), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(18));
    
    hsel2_0_a2_RNIEN1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(15), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(15));
    
    slave_arbiter : COREAHBLITE_SLAVEARBITER_1
      port map(masterAddrInProg(3) => \masterAddrInProg[3]\, 
        masterAddrInProg(2) => \masterAddrInProg[2]\, 
        masterAddrInProg(1) => \masterAddrInProg[1]\, 
        masterAddrInProg(0) => \masterAddrInProg_0\, 
        current_state_0 => current_state_0, xhdl1221_0 => 
        xhdl1221_0, regHMASTLOCK => regHMASTLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        masterRegAddrSel => masterRegAddrSel, SDRCLK_c => 
        SDRCLK_c, MSS_READY => MSS_READY);
    
    hsel2_0_a2_RNIU20O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(6), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(6));
    
    hsel2_0_a2_RNIS00O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(4), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(4));
    
    hwdata10 : CFG4
      generic map(INIT => x"0100")

      port map(A => \masterDataInProg[3]_net_1\, B => 
        \masterDataInProg[2]_net_1\, C => 
        \masterDataInProg[1]_net_1\, D => 
        \masterDataInProg[0]_net_1\, Y => \hwdata10\);
    
    hsel2_0_a2_RNIGQ2T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(26), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(26));
    
    hwdata10_RNILBHG_8 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(22));
    
    hwdata10_RNILBHG_7 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(23));
    
    hsel2_0_a2_RNIAJ1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(11), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(11));
    
    hwdata10_RNILBHG_27 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(3));
    
    hsel2_0_a2_RNIT10O : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(5), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(5));
    
    hsel2_0_a2_RNIBK1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(12), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(12));
    
    hwdata10_RNILBHG_30 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0), B => 
        \hwdata10\, Y => CoreAHBLite_0_AHBmslave10_HWDATA(0));
    
    hsel2_0_a2_RNICL1T : CFG4
      generic map(INIT => x"B800")

      port map(A => regHADDR(13), B => masterRegAddrSel, C => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), D => 
        \hsel2\, Y => CoreAHBLite_0_AHBmslave10_HADDR(13));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_DEFAULTSLAVESM_0 is

    port( DEFSLAVEDATASEL_9      : in    std_logic;
          DEFSLAVEDATASEL_11     : in    std_logic;
          DEFSLAVEDATASEL_10     : in    std_logic;
          defSlaveSMNextState    : out   std_logic;
          SDRCLK_c               : in    std_logic;
          MSS_READY              : in    std_logic;
          defSlaveSMCurrentState : out   std_logic
        );

end COREAHBLITE_DEFAULTSLAVESM_0;

architecture DEF_ARCH of COREAHBLITE_DEFAULTSLAVESM_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal defSlaveSMCurrentState_net_1, VCC_net_1, 
        defSlaveSMNextState_net_1, GND_net_1 : std_logic;

begin 

    defSlaveSMNextState <= defSlaveSMNextState_net_1;
    defSlaveSMCurrentState <= defSlaveSMCurrentState_net_1;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \defSlaveSMNextState\ : CFG4
      generic map(INIT => x"3332")

      port map(A => DEFSLAVEDATASEL_10, B => 
        defSlaveSMCurrentState_net_1, C => DEFSLAVEDATASEL_11, D
         => DEFSLAVEDATASEL_9, Y => defSlaveSMNextState_net_1);
    
    \defSlaveSMCurrentState\ : SLE
      port map(D => defSlaveSMNextState_net_1, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        defSlaveSMCurrentState_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MASTERSTAGE_1_1_0_1024_0 is

    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0);
          regHADDR                                      : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          regHSIZE                                      : out   std_logic_vector(1 downto 0);
          masterAddrInProg_0                            : in    std_logic;
          current_state_0                               : in    std_logic;
          xhdl1292_0                                    : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic;
          xhdl1221_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic;
          N_92                                          : out   std_logic;
          N_91                                          : out   std_logic;
          hready_m_xhdl349                              : out   std_logic;
          masterRegAddrSel                              : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic;
          regHMASTLOCK                                  : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic;
          m0PrevDataSlaveReady                          : out   std_logic;
          SDRCLK_c                                      : in    std_logic;
          MSS_READY                                     : in    std_logic
        );

end COREAHBLITE_MASTERSTAGE_1_1_0_1024_0;

architecture DEF_ARCH of COREAHBLITE_MASTERSTAGE_1_1_0_1024_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_DEFAULTSLAVESM_0
    port( DEFSLAVEDATASEL_9      : in    std_logic := 'U';
          DEFSLAVEDATASEL_11     : in    std_logic := 'U';
          DEFSLAVEDATASEL_10     : in    std_logic := 'U';
          defSlaveSMNextState    : out   std_logic;
          SDRCLK_c               : in    std_logic := 'U';
          MSS_READY              : in    std_logic := 'U';
          defSlaveSMCurrentState : out   std_logic
        );
  end component;

    signal \SDATASELInt[15]_net_1\, VCC_net_1, \SADDRSEL[15]\, 
        \m0PrevDataSlaveReady\, GND_net_1, \SDATASELInt[0]_net_1\, 
        \SADDRSEL[0]\, \SDATASELInt[1]_net_1\, \SADDRSEL[1]\, 
        \SDATASELInt[2]_net_1\, \SADDRSEL[2]\, 
        \SDATASELInt[3]_net_1\, \SADDRSEL[3]\, 
        \SDATASELInt[4]_net_1\, \SADDRSEL[4]\, 
        \SDATASELInt[5]_net_1\, \SADDRSEL[5]\, 
        \SDATASELInt[6]_net_1\, \SADDRSEL[6]\, 
        \SDATASELInt[7]_net_1\, \SADDRSEL[7]\, 
        \SDATASELInt[8]_net_1\, \SADDRSEL[8]\, 
        \SDATASELInt[9]_net_1\, \SADDRSEL[9]\, \xhdl1222_0\, 
        \SDATASELInt_46\, \SDATASELInt[11]_net_1\, \SADDRSEL[11]\, 
        \SDATASELInt[12]_net_1\, \SADDRSEL[12]\, 
        \SDATASELInt[13]_net_1\, \SADDRSEL[13]\, 
        \SDATASELInt[14]_net_1\, \SADDRSEL[14]\, 
        masterAddrClockEnable, \regHADDR[28]_net_1\, 
        \regHADDR[29]_net_1\, \regHADDR[30]_net_1\, 
        \regHADDR[31]_net_1\, \regHWRITE\, \regHTRANS\, 
        masterRegAddrSel_net_1, d_masterRegAddrSel, \HRESP_0_am\, 
        \hready_m_xhdl349\, un1_hready_m_xhdl339_i, 
        \M0GATEDHADDR[30]\, \M0GATEDHADDR[29]\, G_11_1, 
        \M0GATEDHADDR[28]\, \xhdl1221_0\, \M0GATEDHADDR[31]\, 
        \SADDRSEL_0_a2_0_0[2]_net_1\, \N_92\, 
        \d_masterRegAddrSel_0_a2_0\, \DEFSLAVEDATASEL_10\, 
        \DEFSLAVEDATASEL_9\, \DEFSLAVEDATASEL_8\, N_3059, N_3060, 
        N_66, N_67, N_150, N_139, \masterAddrClockEnable_0_a2_1\, 
        \DEFSLAVEDATASEL_11\, N_3062, N_3042, N_17, N_3043, N_19, 
        N_3045, N_3048, \un1_hready_m_xhdl339_0_0_1_tz\, 
        \un1_hready_m_xhdl339_0_0_1\, defSlaveSMCurrentState, 
        defSlaveSMNextState, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY\, 
        \masterAddrClockEnable_0_a2_2\, 
        \d_masterRegAddrSel_0_a2_1\ : std_logic;

    for all : COREAHBLITE_DEFAULTSLAVESM_0
	Use entity work.COREAHBLITE_DEFAULTSLAVESM_0(DEF_ARCH);
begin 

    xhdl1221_0 <= \xhdl1221_0\;
    xhdl1222_0 <= \xhdl1222_0\;
    top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY <= 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY\;
    N_92 <= \N_92\;
    hready_m_xhdl349 <= \hready_m_xhdl349\;
    masterRegAddrSel <= masterRegAddrSel_net_1;
    m0PrevDataSlaveReady <= \m0PrevDataSlaveReady\;

    \regHADDR[21]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(21));
    
    \PREGATEDHADDR[31]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31), C => 
        \regHADDR[31]_net_1\, Y => \M0GATEDHADDR[31]\);
    
    \regHADDR[15]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(15));
    
    \regHADDR[30]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \regHADDR[30]_net_1\);
    
    DEFSLAVEDATASEL_10 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[12]_net_1\, C => \SDATASELInt[11]_net_1\, D
         => \SDATASELInt[9]_net_1\, Y => \DEFSLAVEDATASEL_10\);
    
    \regHADDR[7]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(7));
    
    un1_hready_m_xhdl339_0_o2 : CFG3
      generic map(INIT => x"16")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[13]_net_1\, C => \SDATASELInt[9]_net_1\, Y
         => N_3042);
    
    \SADDRSEL_0_a2[6]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \M0GATEDHADDR[28]\, B => N_150, C => 
        \M0GATEDHADDR[31]\, Y => \SADDRSEL[6]\);
    
    \SADDRSEL_0_a2[0]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[0]\);
    
    \PREGATEDHADDR[30]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30), C => 
        \regHADDR[30]_net_1\, Y => \M0GATEDHADDR[30]\);
    
    un1_hready_m_xhdl339_0_0_1 : CFG4
      generic map(INIT => x"0800")

      port map(A => N_3059, B => \un1_hready_m_xhdl339_0_0_1_tz\, 
        C => \xhdl1222_0\, D => N_67, Y => 
        \un1_hready_m_xhdl339_0_0_1\);
    
    \SADDRSEL_0_a2_0[14]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \M0GATEDHADDR[29]\, B => \M0GATEDHADDR[30]\, 
        C => \N_92\, Y => N_150);
    
    regHTRANS_RNI9J371 : CFG4
      generic map(INIT => x"3F77")

      port map(A => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, 
        B => \M0GATEDHADDR[31]\, C => \regHTRANS\, D => 
        masterRegAddrSel_net_1, Y => G_11_1);
    
    \regHADDR[9]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(9));
    
    \SADDRSEL_0_a2[3]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \M0GATEDHADDR[31]\, B => \M0GATEDHADDR[28]\, 
        C => \N_92\, D => \SADDRSEL_0_a2_0_0[2]_net_1\, Y => 
        \SADDRSEL[3]\);
    
    \masterRegAddrSel\ : SLE
      port map(D => d_masterRegAddrSel, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        masterRegAddrSel_net_1);
    
    masterAddrClockEnable_0_a2_2 : CFG3
      generic map(INIT => x"80")

      port map(A => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, 
        B => \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY\, C => 
        \masterAddrClockEnable_0_a2_1\, Y => 
        \masterAddrClockEnable_0_a2_2\);
    
    \SADDRSEL_0_a2[15]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \M0GATEDHADDR[28]\, B => N_150, C => 
        \M0GATEDHADDR[31]\, Y => \SADDRSEL[15]\);
    
    regHTRANS : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => 
        masterAddrClockEnable, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \regHTRANS\);
    
    \SADDRSEL_0_a2_0_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \M0GATEDHADDR[30]\, B => \M0GATEDHADDR[29]\, 
        Y => \SADDRSEL_0_a2_0_0[2]_net_1\);
    
    GATEDHTRANS_i_m2 : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, C => 
        \regHTRANS\, Y => \N_92\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un1_hready_m_xhdl339_0_a2_13 : CFG3
      generic map(INIT => x"01")

      port map(A => \SDATASELInt[14]_net_1\, B => 
        \SDATASELInt[13]_net_1\, C => \SDATASELInt[9]_net_1\, Y
         => N_67);
    
    \SADDRSEL_0_a2[12]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[12]\);
    
    \SADDRSEL_0_a2[4]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[4]\);
    
    \regHADDR[29]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \regHADDR[29]_net_1\);
    
    hready_m_xhdl349_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => \xhdl1222_0\, B => N_67, C => N_3059, D => 
        N_3062, Y => \hready_m_xhdl349\);
    
    d_masterRegAddrSel_0_a2_0 : CFG3
      generic map(INIT => x"40")

      port map(A => \M0GATEDHADDR[28]\, B => 
        \SADDRSEL_0_a2_0_0[2]_net_1\, C => \M0GATEDHADDR[31]\, Y
         => \d_masterRegAddrSel_0_a2_0\);
    
    \regHADDR[24]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(24));
    
    \SADDRSEL_0_a2[14]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \M0GATEDHADDR[28]\, B => N_150, C => 
        \M0GATEDHADDR[31]\, Y => \SADDRSEL[14]\);
    
    \regHADDR[28]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \regHADDR[28]_net_1\);
    
    SDATASELInt_46 : CFG3
      generic map(INIT => x"AC")

      port map(A => \xhdl1221_0\, B => \xhdl1222_0\, C => 
        \m0PrevDataSlaveReady\, Y => \SDATASELInt_46\);
    
    \regHADDR[31]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \regHADDR[31]_net_1\);
    
    \regHADDR[10]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(10));
    
    \SADDRSEL_0_a2[8]\ : CFG4
      generic map(INIT => x"0400")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[8]\);
    
    \regHADDR[13]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(13));
    
    \regHADDR[12]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(12));
    
    HRESP_0_am : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \DEFSLAVEDATASEL_10\, B => 
        defSlaveSMCurrentState, C => \DEFSLAVEDATASEL_11\, D => 
        \DEFSLAVEDATASEL_9\, Y => \HRESP_0_am\);
    
    \regHADDR[5]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(5));
    
    \SDATASELInt[4]\ : SLE
      port map(D => \SADDRSEL[4]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[4]_net_1\);
    
    \regHADDR[2]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(2));
    
    \SDATASELInt[15]\ : SLE
      port map(D => \SADDRSEL[15]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[15]_net_1\);
    
    \PREGATEDHADDR[28]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28), C => 
        \regHADDR[28]_net_1\, Y => \M0GATEDHADDR[28]\);
    
    \SDATASELInt[14]\ : SLE
      port map(D => \SADDRSEL[14]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[14]_net_1\);
    
    GATEDHWRITE_i_m2 : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, C => 
        \regHWRITE\, Y => N_91);
    
    \SDATASELInt[2]\ : SLE
      port map(D => \SADDRSEL[2]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[2]_net_1\);
    
    \regHADDR[8]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(8));
    
    \regHADDR[25]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(25));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    hready_m_xhdl349_0_a2_0 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[12]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \SDATASELInt[1]_net_1\, D
         => \SDATASELInt[0]_net_1\, Y => N_3059);
    
    \regHADDR[17]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(17));
    
    un1_hready_m_xhdl339_0_a2_12 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[11]_net_1\, C => \SDATASELInt[8]_net_1\, D
         => \SDATASELInt[7]_net_1\, Y => N_66);
    
    \SADDRSEL_0_a2[7]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \M0GATEDHADDR[28]\, B => N_150, C => 
        \M0GATEDHADDR[31]\, Y => \SADDRSEL[7]\);
    
    \regHADDR[6]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(6));
    
    \regHADDR[16]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(16));
    
    DEFSLAVEDATASEL_9 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \SDATASELInt[13]_net_1\, B => 
        \SDATASELInt[8]_net_1\, C => \SDATASELInt[7]_net_1\, D
         => \SDATASELInt[6]_net_1\, Y => \DEFSLAVEDATASEL_9\);
    
    \SDATASELInt[13]\ : SLE
      port map(D => \SADDRSEL[13]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[13]_net_1\);
    
    \SADDRSEL_0_a2[11]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \M0GATEDHADDR[31]\, B => \M0GATEDHADDR[28]\, 
        C => \N_92\, D => \SADDRSEL_0_a2_0_0[2]_net_1\, Y => 
        \SADDRSEL[11]\);
    
    un1_hready_m_xhdl339_0_o2_1 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[6]_net_1\, B => 
        \SDATASELInt[5]_net_1\, C => \SDATASELInt[4]_net_1\, D
         => \SDATASELInt[3]_net_1\, Y => N_3043);
    
    regHWRITE : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \regHWRITE\);
    
    \regHSIZE[1]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHSIZE(1));
    
    \regHMASTLOCK\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHMASTLOCK);
    
    \SDATASELInt[9]\ : SLE
      port map(D => \SADDRSEL[9]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[9]_net_1\);
    
    \SDATASELInt[1]\ : SLE
      port map(D => \SADDRSEL[1]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[1]_net_1\);
    
    \SDATASELInt[12]\ : SLE
      port map(D => \SADDRSEL[12]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[12]_net_1\);
    
    \SDATASELInt[0]\ : SLE
      port map(D => \SADDRSEL[0]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[0]_net_1\);
    
    \regHADDR[11]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(11));
    
    \regHADDR[0]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(0));
    
    \SDATASELInt[5]\ : SLE
      port map(D => \SADDRSEL[5]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[5]_net_1\);
    
    \PREGATEDHADDR_RNIOOFI2[29]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \M0GATEDHADDR[30]\, B => \M0GATEDHADDR[29]\, 
        C => G_11_1, D => \M0GATEDHADDR[28]\, Y => \xhdl1221_0\);
    
    masterAddrClockEnable_0_a2_1 : CFG4
      generic map(INIT => x"0020")

      port map(A => \M0GATEDHADDR[31]\, B => 
        masterRegAddrSel_net_1, C => \SADDRSEL_0_a2_0_0[2]_net_1\, 
        D => \M0GATEDHADDR[28]\, Y => 
        \masterAddrClockEnable_0_a2_1\);
    
    HRESP_u : CFG3
      generic map(INIT => x"20")

      port map(A => \HRESP_0_am\, B => \hready_m_xhdl349\, C => 
        un1_hready_m_xhdl339_i, Y => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0);
    
    \regHADDR[3]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(3));
    
    \SADDRSEL_0_a2[5]\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[5]\);
    
    un1_hready_m_xhdl339_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => \xhdl1222_0\, B => N_19, C => N_67, D => 
        N_3062, Y => N_3045);
    
    \SDATASELInt[3]\ : SLE
      port map(D => \SADDRSEL[3]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[3]_net_1\);
    
    d_masterRegAddrSel_0_a2_1 : CFG4
      generic map(INIT => x"E0C0")

      port map(A => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, 
        B => masterRegAddrSel_net_1, C => 
        \d_masterRegAddrSel_0_a2_0\, D => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY\, Y => 
        \d_masterRegAddrSel_0_a2_1\);
    
    un1_hready_m_xhdl339_0_a2_2 : CFG4
      generic map(INIT => x"4000")

      port map(A => \xhdl1222_0\, B => N_3042, C => N_3059, D => 
        N_3062, Y => N_3048);
    
    un1_hready_m_xhdl339_0_0 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => N_3048, B => \un1_hready_m_xhdl339_0_0_1\, C
         => \hready_m_xhdl349\, D => N_3045, Y => 
        un1_hready_m_xhdl339_i);
    
    un1_hready_m_xhdl339_0_0_1_tz : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_3043, B => N_17, C => N_3060, D => N_66, Y
         => \un1_hready_m_xhdl339_0_0_1_tz\);
    
    \regHADDR[20]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(20));
    
    un1_hready_m_xhdl339_0_a2_11 : CFG4
      generic map(INIT => x"0001")

      port map(A => \SDATASELInt[6]_net_1\, B => 
        \SDATASELInt[5]_net_1\, C => \SDATASELInt[4]_net_1\, D
         => \SDATASELInt[3]_net_1\, Y => N_3060);
    
    \SADDRSEL_0_a2_2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \N_92\, B => \M0GATEDHADDR[29]\, Y => N_139);
    
    \regHADDR[23]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(23));
    
    \regHADDR[1]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(1));
    
    \regHADDR[22]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(22));
    
    \SDATASELInt[7]\ : SLE
      port map(D => \SADDRSEL[7]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[7]_net_1\);
    
    \regHSIZE[0]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHSIZE(0));
    
    un1_hready_m_xhdl339_0_a2_14 : CFG2
      generic map(INIT => x"8")

      port map(A => N_66, B => N_3060, Y => N_3062);
    
    \SADDRSEL_0_a2[1]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[1]\);
    
    \SADDRSEL_0_a2[13]\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[13]\);
    
    DEFSLAVEDATASEL_8 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \SDATASELInt[5]_net_1\, B => 
        \SDATASELInt[4]_net_1\, C => \SDATASELInt[3]_net_1\, D
         => \SDATASELInt[2]_net_1\, Y => \DEFSLAVEDATASEL_8\);
    
    \SDATASELInt[6]\ : SLE
      port map(D => \SADDRSEL[6]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[6]_net_1\);
    
    \PREGATEDHADDR[29]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => masterRegAddrSel_net_1, B => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29), C => 
        \regHADDR[29]_net_1\, Y => \M0GATEDHADDR[29]\);
    
    PREVDATASLAVEREADY_u : CFG4
      generic map(INIT => x"B3F7")

      port map(A => \hready_m_xhdl349\, B => 
        un1_hready_m_xhdl339_i, C => current_state_0, D => 
        defSlaveSMNextState, Y => \m0PrevDataSlaveReady\);
    
    \regHADDR[19]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(19));
    
    \regHADDR[14]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(14));
    
    HREADY_M_u : CFG4
      generic map(INIT => x"B3F7")

      port map(A => \hready_m_xhdl349\, B => 
        un1_hready_m_xhdl339_i, C => xhdl1292_0, D => 
        defSlaveSMNextState, Y => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY\);
    
    d_masterRegAddrSel_0_a2 : CFG4
      generic map(INIT => x"2A00")

      port map(A => \xhdl1221_0\, B => current_state_0, C => 
        masterAddrInProg_0, D => \d_masterRegAddrSel_0_a2_1\, Y
         => d_masterRegAddrSel);
    
    \SADDRSEL_0_a2[2]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \M0GATEDHADDR[31]\, B => \M0GATEDHADDR[28]\, 
        C => \N_92\, D => \SADDRSEL_0_a2_0_0[2]_net_1\, Y => 
        \SADDRSEL[2]\);
    
    \regHADDR[27]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(27));
    
    un1_hready_m_xhdl339_0_o2_0 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[11]_net_1\, C => \SDATASELInt[8]_net_1\, D
         => \SDATASELInt[7]_net_1\, Y => N_17);
    
    \regHADDR[18]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(18));
    
    \SDATASELInt[11]\ : SLE
      port map(D => \SADDRSEL[11]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[11]_net_1\);
    
    DEFSLAVEDATASEL_11 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \SDATASELInt[15]_net_1\, B => 
        \SDATASELInt[1]_net_1\, C => \SDATASELInt[0]_net_1\, D
         => \DEFSLAVEDATASEL_8\, Y => \DEFSLAVEDATASEL_11\);
    
    un1_hready_m_xhdl339_0_o2_2 : CFG4
      generic map(INIT => x"0116")

      port map(A => \SDATASELInt[12]_net_1\, B => 
        \SDATASELInt[2]_net_1\, C => \SDATASELInt[1]_net_1\, D
         => \SDATASELInt[0]_net_1\, Y => N_19);
    
    \SDATASELInt[8]\ : SLE
      port map(D => \SADDRSEL[8]\, CLK => SDRCLK_c, EN => 
        \m0PrevDataSlaveReady\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \SDATASELInt[8]_net_1\);
    
    \regHADDR[4]\ : SLE
      port map(D => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), 
        CLK => SDRCLK_c, EN => masterAddrClockEnable, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => regHADDR(4));
    
    \regHADDR[26]\ : SLE
      port map(D => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), CLK => 
        SDRCLK_c, EN => masterAddrClockEnable, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => regHADDR(26));
    
    \SDATASELInt[10]\ : SLE
      port map(D => \SDATASELInt_46\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \xhdl1222_0\);
    
    masterAddrClockEnable_0_a2 : CFG4
      generic map(INIT => x"2A00")

      port map(A => \xhdl1221_0\, B => current_state_0, C => 
        masterAddrInProg_0, D => \masterAddrClockEnable_0_a2_2\, 
        Y => masterAddrClockEnable);
    
    \SADDRSEL_0_a2[9]\ : CFG4
      generic map(INIT => x"0800")

      port map(A => \M0GATEDHADDR[28]\, B => N_139, C => 
        \M0GATEDHADDR[30]\, D => \M0GATEDHADDR[31]\, Y => 
        \SADDRSEL[9]\);
    
    default_slave_sm : COREAHBLITE_DEFAULTSLAVESM_0
      port map(DEFSLAVEDATASEL_9 => \DEFSLAVEDATASEL_9\, 
        DEFSLAVEDATASEL_11 => \DEFSLAVEDATASEL_11\, 
        DEFSLAVEDATASEL_10 => \DEFSLAVEDATASEL_10\, 
        defSlaveSMNextState => defSlaveSMNextState, SDRCLK_c => 
        SDRCLK_c, MSS_READY => MSS_READY, defSlaveSMCurrentState
         => defSlaveSMCurrentState);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity COREAHBLITE_MATRIX4X16 is

    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA              : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE               : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HADDR               : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0);
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic;
          current_state_0                               : in    std_logic;
          masterAddrInProg_0                            : out   std_logic;
          hsel2_0_a2_1                                  : out   std_logic;
          hsel2                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE              : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK           : out   std_logic;
          MSS_READY                                     : in    std_logic;
          SDRCLK_c                                      : in    std_logic;
          m0PrevDataSlaveReady                          : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic;
          hready_m_xhdl349                              : out   std_logic;
          N_91                                          : out   std_logic;
          N_92                                          : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic
        );

end COREAHBLITE_MATRIX4X16;

architecture DEF_ARCH of COREAHBLITE_MATRIX4X16 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_SLAVESTAGE_0
    port( CoreAHBLite_0_AHBmslave10_HADDR             : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR  : in    std_logic_vector(27 downto 0) := (others => 'U');
          regHADDR                                    : in    std_logic_vector(27 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HSIZE             : out   std_logic_vector(1 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE  : in    std_logic_vector(1 downto 0) := (others => 'U');
          regHSIZE                                    : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HWDATA            : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA : in    std_logic_vector(31 downto 0) := (others => 'U');
          xhdl1221_0                                  : in    std_logic := 'U';
          masterAddrInProg_0                          : out   std_logic;
          xhdl1292_0                                  : out   std_logic;
          xhdl1222_0                                  : in    std_logic := 'U';
          current_state_0                             : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave10_HMASTLOCK         : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK  : in    std_logic := 'U';
          masterRegAddrSel                            : in    std_logic := 'U';
          regHMASTLOCK                                : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave10_HWRITE            : out   std_logic;
          N_91                                        : in    std_logic := 'U';
          hsel2                                       : out   std_logic;
          hsel2_0_a2_1                                : out   std_logic;
          SDRCLK_c                                    : in    std_logic := 'U';
          MSS_READY                                   : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MASTERSTAGE_1_1_0_1024_0
    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0) := (others => 'U');
          regHADDR                                      : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          regHSIZE                                      : out   std_logic_vector(1 downto 0);
          masterAddrInProg_0                            : in    std_logic := 'U';
          current_state_0                               : in    std_logic := 'U';
          xhdl1292_0                                    : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic := 'U';
          xhdl1221_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic;
          N_92                                          : out   std_logic;
          N_91                                          : out   std_logic;
          hready_m_xhdl349                              : out   std_logic;
          masterRegAddrSel                              : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic := 'U';
          regHMASTLOCK                                  : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          m0PrevDataSlaveReady                          : out   std_logic;
          SDRCLK_c                                      : in    std_logic := 'U';
          MSS_READY                                     : in    std_logic := 'U'
        );
  end component;

    signal \masterAddrInProg_0\, \xhdl1292[0]\, \xhdl1221[10]\, 
        \regHADDR[0]\, \regHADDR[1]\, \regHADDR[2]\, 
        \regHADDR[3]\, \regHADDR[4]\, \regHADDR[5]\, 
        \regHADDR[6]\, \regHADDR[7]\, \regHADDR[8]\, 
        \regHADDR[9]\, \regHADDR[10]\, \regHADDR[11]\, 
        \regHADDR[12]\, \regHADDR[13]\, \regHADDR[14]\, 
        \regHADDR[15]\, \regHADDR[16]\, \regHADDR[17]\, 
        \regHADDR[18]\, \regHADDR[19]\, \regHADDR[20]\, 
        \regHADDR[21]\, \regHADDR[22]\, \regHADDR[23]\, 
        \regHADDR[24]\, \regHADDR[25]\, \regHADDR[26]\, 
        \regHADDR[27]\, \regHSIZE[0]\, \regHSIZE[1]\, 
        \xhdl1222_0\, \N_91\, masterRegAddrSel, regHMASTLOCK, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_SLAVESTAGE_0
	Use entity work.COREAHBLITE_SLAVESTAGE_0(DEF_ARCH);
    for all : COREAHBLITE_MASTERSTAGE_1_1_0_1024_0
	Use entity work.COREAHBLITE_MASTERSTAGE_1_1_0_1024_0(DEF_ARCH);
begin 

    xhdl1222_0 <= \xhdl1222_0\;
    masterAddrInProg_0 <= \masterAddrInProg_0\;
    N_91 <= \N_91\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    slavestage_10 : COREAHBLITE_SLAVESTAGE_0
      port map(CoreAHBLite_0_AHBmslave10_HADDR(27) => 
        CoreAHBLite_0_AHBmslave10_HADDR(27), 
        CoreAHBLite_0_AHBmslave10_HADDR(26) => 
        CoreAHBLite_0_AHBmslave10_HADDR(26), 
        CoreAHBLite_0_AHBmslave10_HADDR(25) => 
        CoreAHBLite_0_AHBmslave10_HADDR(25), 
        CoreAHBLite_0_AHBmslave10_HADDR(24) => 
        CoreAHBLite_0_AHBmslave10_HADDR(24), 
        CoreAHBLite_0_AHBmslave10_HADDR(23) => 
        CoreAHBLite_0_AHBmslave10_HADDR(23), 
        CoreAHBLite_0_AHBmslave10_HADDR(22) => 
        CoreAHBLite_0_AHBmslave10_HADDR(22), 
        CoreAHBLite_0_AHBmslave10_HADDR(21) => 
        CoreAHBLite_0_AHBmslave10_HADDR(21), 
        CoreAHBLite_0_AHBmslave10_HADDR(20) => 
        CoreAHBLite_0_AHBmslave10_HADDR(20), 
        CoreAHBLite_0_AHBmslave10_HADDR(19) => 
        CoreAHBLite_0_AHBmslave10_HADDR(19), 
        CoreAHBLite_0_AHBmslave10_HADDR(18) => 
        CoreAHBLite_0_AHBmslave10_HADDR(18), 
        CoreAHBLite_0_AHBmslave10_HADDR(17) => 
        CoreAHBLite_0_AHBmslave10_HADDR(17), 
        CoreAHBLite_0_AHBmslave10_HADDR(16) => 
        CoreAHBLite_0_AHBmslave10_HADDR(16), 
        CoreAHBLite_0_AHBmslave10_HADDR(15) => 
        CoreAHBLite_0_AHBmslave10_HADDR(15), 
        CoreAHBLite_0_AHBmslave10_HADDR(14) => 
        CoreAHBLite_0_AHBmslave10_HADDR(14), 
        CoreAHBLite_0_AHBmslave10_HADDR(13) => 
        CoreAHBLite_0_AHBmslave10_HADDR(13), 
        CoreAHBLite_0_AHBmslave10_HADDR(12) => 
        CoreAHBLite_0_AHBmslave10_HADDR(12), 
        CoreAHBLite_0_AHBmslave10_HADDR(11) => 
        CoreAHBLite_0_AHBmslave10_HADDR(11), 
        CoreAHBLite_0_AHBmslave10_HADDR(10) => 
        CoreAHBLite_0_AHBmslave10_HADDR(10), 
        CoreAHBLite_0_AHBmslave10_HADDR(9) => 
        CoreAHBLite_0_AHBmslave10_HADDR(9), 
        CoreAHBLite_0_AHBmslave10_HADDR(8) => 
        CoreAHBLite_0_AHBmslave10_HADDR(8), 
        CoreAHBLite_0_AHBmslave10_HADDR(7) => 
        CoreAHBLite_0_AHBmslave10_HADDR(7), 
        CoreAHBLite_0_AHBmslave10_HADDR(6) => 
        CoreAHBLite_0_AHBmslave10_HADDR(6), 
        CoreAHBLite_0_AHBmslave10_HADDR(5) => 
        CoreAHBLite_0_AHBmslave10_HADDR(5), 
        CoreAHBLite_0_AHBmslave10_HADDR(4) => 
        CoreAHBLite_0_AHBmslave10_HADDR(4), 
        CoreAHBLite_0_AHBmslave10_HADDR(3) => 
        CoreAHBLite_0_AHBmslave10_HADDR(3), 
        CoreAHBLite_0_AHBmslave10_HADDR(2) => 
        CoreAHBLite_0_AHBmslave10_HADDR(2), 
        CoreAHBLite_0_AHBmslave10_HADDR(1) => 
        CoreAHBLite_0_AHBmslave10_HADDR(1), 
        CoreAHBLite_0_AHBmslave10_HADDR(0) => 
        CoreAHBLite_0_AHBmslave10_HADDR(0), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), 
        regHADDR(27) => \regHADDR[27]\, regHADDR(26) => 
        \regHADDR[26]\, regHADDR(25) => \regHADDR[25]\, 
        regHADDR(24) => \regHADDR[24]\, regHADDR(23) => 
        \regHADDR[23]\, regHADDR(22) => \regHADDR[22]\, 
        regHADDR(21) => \regHADDR[21]\, regHADDR(20) => 
        \regHADDR[20]\, regHADDR(19) => \regHADDR[19]\, 
        regHADDR(18) => \regHADDR[18]\, regHADDR(17) => 
        \regHADDR[17]\, regHADDR(16) => \regHADDR[16]\, 
        regHADDR(15) => \regHADDR[15]\, regHADDR(14) => 
        \regHADDR[14]\, regHADDR(13) => \regHADDR[13]\, 
        regHADDR(12) => \regHADDR[12]\, regHADDR(11) => 
        \regHADDR[11]\, regHADDR(10) => \regHADDR[10]\, 
        regHADDR(9) => \regHADDR[9]\, regHADDR(8) => 
        \regHADDR[8]\, regHADDR(7) => \regHADDR[7]\, regHADDR(6)
         => \regHADDR[6]\, regHADDR(5) => \regHADDR[5]\, 
        regHADDR(4) => \regHADDR[4]\, regHADDR(3) => 
        \regHADDR[3]\, regHADDR(2) => \regHADDR[2]\, regHADDR(1)
         => \regHADDR[1]\, regHADDR(0) => \regHADDR[0]\, 
        CoreAHBLite_0_AHBmslave10_HSIZE(1) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(1), 
        CoreAHBLite_0_AHBmslave10_HSIZE(0) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(0), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), 
        regHSIZE(1) => \regHSIZE[1]\, regHSIZE(0) => 
        \regHSIZE[0]\, CoreAHBLite_0_AHBmslave10_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(31), 
        CoreAHBLite_0_AHBmslave10_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(30), 
        CoreAHBLite_0_AHBmslave10_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(29), 
        CoreAHBLite_0_AHBmslave10_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(28), 
        CoreAHBLite_0_AHBmslave10_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(27), 
        CoreAHBLite_0_AHBmslave10_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(26), 
        CoreAHBLite_0_AHBmslave10_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(25), 
        CoreAHBLite_0_AHBmslave10_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(24), 
        CoreAHBLite_0_AHBmslave10_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(23), 
        CoreAHBLite_0_AHBmslave10_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(22), 
        CoreAHBLite_0_AHBmslave10_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(21), 
        CoreAHBLite_0_AHBmslave10_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(20), 
        CoreAHBLite_0_AHBmslave10_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(19), 
        CoreAHBLite_0_AHBmslave10_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(18), 
        CoreAHBLite_0_AHBmslave10_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(17), 
        CoreAHBLite_0_AHBmslave10_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(16), 
        CoreAHBLite_0_AHBmslave10_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(15), 
        CoreAHBLite_0_AHBmslave10_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(14), 
        CoreAHBLite_0_AHBmslave10_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(13), 
        CoreAHBLite_0_AHBmslave10_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(12), 
        CoreAHBLite_0_AHBmslave10_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(11), 
        CoreAHBLite_0_AHBmslave10_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(10), 
        CoreAHBLite_0_AHBmslave10_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(9), 
        CoreAHBLite_0_AHBmslave10_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(8), 
        CoreAHBLite_0_AHBmslave10_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(7), 
        CoreAHBLite_0_AHBmslave10_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(6), 
        CoreAHBLite_0_AHBmslave10_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(5), 
        CoreAHBLite_0_AHBmslave10_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(4), 
        CoreAHBLite_0_AHBmslave10_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(3), 
        CoreAHBLite_0_AHBmslave10_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(2), 
        CoreAHBLite_0_AHBmslave10_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(1), 
        CoreAHBLite_0_AHBmslave10_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(0), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0), 
        xhdl1221_0 => \xhdl1221[10]\, masterAddrInProg_0 => 
        \masterAddrInProg_0\, xhdl1292_0 => \xhdl1292[0]\, 
        xhdl1222_0 => \xhdl1222_0\, current_state_0 => 
        current_state_0, CoreAHBLite_0_AHBmslave10_HMASTLOCK => 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        masterRegAddrSel => masterRegAddrSel, regHMASTLOCK => 
        regHMASTLOCK, CoreAHBLite_0_AHBmslave10_HWRITE => 
        CoreAHBLite_0_AHBmslave10_HWRITE, N_91 => \N_91\, hsel2
         => hsel2, hsel2_0_a2_1 => hsel2_0_a2_1, SDRCLK_c => 
        SDRCLK_c, MSS_READY => MSS_READY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    masterstage_0 : COREAHBLITE_MASTERSTAGE_1_1_0_1024_0
      port map(top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), 
        regHADDR(27) => \regHADDR[27]\, regHADDR(26) => 
        \regHADDR[26]\, regHADDR(25) => \regHADDR[25]\, 
        regHADDR(24) => \regHADDR[24]\, regHADDR(23) => 
        \regHADDR[23]\, regHADDR(22) => \regHADDR[22]\, 
        regHADDR(21) => \regHADDR[21]\, regHADDR(20) => 
        \regHADDR[20]\, regHADDR(19) => \regHADDR[19]\, 
        regHADDR(18) => \regHADDR[18]\, regHADDR(17) => 
        \regHADDR[17]\, regHADDR(16) => \regHADDR[16]\, 
        regHADDR(15) => \regHADDR[15]\, regHADDR(14) => 
        \regHADDR[14]\, regHADDR(13) => \regHADDR[13]\, 
        regHADDR(12) => \regHADDR[12]\, regHADDR(11) => 
        \regHADDR[11]\, regHADDR(10) => \regHADDR[10]\, 
        regHADDR(9) => \regHADDR[9]\, regHADDR(8) => 
        \regHADDR[8]\, regHADDR(7) => \regHADDR[7]\, regHADDR(6)
         => \regHADDR[6]\, regHADDR(5) => \regHADDR[5]\, 
        regHADDR(4) => \regHADDR[4]\, regHADDR(3) => 
        \regHADDR[3]\, regHADDR(2) => \regHADDR[2]\, regHADDR(1)
         => \regHADDR[1]\, regHADDR(0) => \regHADDR[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), 
        regHSIZE(1) => \regHSIZE[1]\, regHSIZE(0) => 
        \regHSIZE[0]\, masterAddrInProg_0 => \masterAddrInProg_0\, 
        current_state_0 => current_state_0, xhdl1292_0 => 
        \xhdl1292[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, xhdl1221_0
         => \xhdl1221[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0 => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0, xhdl1222_0
         => \xhdl1222_0\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY, N_92 => N_92, 
        N_91 => \N_91\, hready_m_xhdl349 => hready_m_xhdl349, 
        masterRegAddrSel => masterRegAddrSel, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, regHMASTLOCK
         => regHMASTLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        m0PrevDataSlaveReady => m0PrevDataSlaveReady, SDRCLK_c
         => SDRCLK_c, MSS_READY => MSS_READY);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLite is

    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HADDR               : out   std_logic_vector(27 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE               : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA              : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0);
          masterAddrInProg_0                            : out   std_logic;
          current_state_0                               : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic;
          N_92                                          : out   std_logic;
          N_91                                          : out   std_logic;
          hready_m_xhdl349                              : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic;
          m0PrevDataSlaveReady                          : out   std_logic;
          SDRCLK_c                                      : in    std_logic;
          MSS_READY                                     : in    std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK           : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE              : out   std_logic;
          hsel2                                         : out   std_logic;
          hsel2_0_a2_1                                  : out   std_logic
        );

end CoreAHBLite;

architecture DEF_ARCH of CoreAHBLite is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component COREAHBLITE_MATRIX4X16
    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HWDATA              : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE               : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HADDR               : out   std_logic_vector(27 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0) := (others => 'U');
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic := 'U';
          current_state_0                               : in    std_logic := 'U';
          masterAddrInProg_0                            : out   std_logic;
          hsel2_0_a2_1                                  : out   std_logic;
          hsel2                                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE              : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK           : out   std_logic;
          MSS_READY                                     : in    std_logic := 'U';
          SDRCLK_c                                      : in    std_logic := 'U';
          m0PrevDataSlaveReady                          : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic := 'U';
          hready_m_xhdl349                              : out   std_logic;
          N_91                                          : out   std_logic;
          N_92                                          : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : COREAHBLITE_MATRIX4X16
	Use entity work.COREAHBLITE_MATRIX4X16(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    matrix4x16 : COREAHBLITE_MATRIX4X16
      port map(top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31)
         => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0), 
        CoreAHBLite_0_AHBmslave10_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(31), 
        CoreAHBLite_0_AHBmslave10_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(30), 
        CoreAHBLite_0_AHBmslave10_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(29), 
        CoreAHBLite_0_AHBmslave10_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(28), 
        CoreAHBLite_0_AHBmslave10_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(27), 
        CoreAHBLite_0_AHBmslave10_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(26), 
        CoreAHBLite_0_AHBmslave10_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(25), 
        CoreAHBLite_0_AHBmslave10_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(24), 
        CoreAHBLite_0_AHBmslave10_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(23), 
        CoreAHBLite_0_AHBmslave10_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(22), 
        CoreAHBLite_0_AHBmslave10_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(21), 
        CoreAHBLite_0_AHBmslave10_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(20), 
        CoreAHBLite_0_AHBmslave10_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(19), 
        CoreAHBLite_0_AHBmslave10_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(18), 
        CoreAHBLite_0_AHBmslave10_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(17), 
        CoreAHBLite_0_AHBmslave10_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(16), 
        CoreAHBLite_0_AHBmslave10_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(15), 
        CoreAHBLite_0_AHBmslave10_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(14), 
        CoreAHBLite_0_AHBmslave10_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(13), 
        CoreAHBLite_0_AHBmslave10_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(12), 
        CoreAHBLite_0_AHBmslave10_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(11), 
        CoreAHBLite_0_AHBmslave10_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(10), 
        CoreAHBLite_0_AHBmslave10_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(9), 
        CoreAHBLite_0_AHBmslave10_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(8), 
        CoreAHBLite_0_AHBmslave10_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(7), 
        CoreAHBLite_0_AHBmslave10_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(6), 
        CoreAHBLite_0_AHBmslave10_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(5), 
        CoreAHBLite_0_AHBmslave10_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(4), 
        CoreAHBLite_0_AHBmslave10_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(3), 
        CoreAHBLite_0_AHBmslave10_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(2), 
        CoreAHBLite_0_AHBmslave10_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(1), 
        CoreAHBLite_0_AHBmslave10_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(0), 
        CoreAHBLite_0_AHBmslave10_HSIZE(1) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(1), 
        CoreAHBLite_0_AHBmslave10_HSIZE(0) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(0), 
        CoreAHBLite_0_AHBmslave10_HADDR(27) => 
        CoreAHBLite_0_AHBmslave10_HADDR(27), 
        CoreAHBLite_0_AHBmslave10_HADDR(26) => 
        CoreAHBLite_0_AHBmslave10_HADDR(26), 
        CoreAHBLite_0_AHBmslave10_HADDR(25) => 
        CoreAHBLite_0_AHBmslave10_HADDR(25), 
        CoreAHBLite_0_AHBmslave10_HADDR(24) => 
        CoreAHBLite_0_AHBmslave10_HADDR(24), 
        CoreAHBLite_0_AHBmslave10_HADDR(23) => 
        CoreAHBLite_0_AHBmslave10_HADDR(23), 
        CoreAHBLite_0_AHBmslave10_HADDR(22) => 
        CoreAHBLite_0_AHBmslave10_HADDR(22), 
        CoreAHBLite_0_AHBmslave10_HADDR(21) => 
        CoreAHBLite_0_AHBmslave10_HADDR(21), 
        CoreAHBLite_0_AHBmslave10_HADDR(20) => 
        CoreAHBLite_0_AHBmslave10_HADDR(20), 
        CoreAHBLite_0_AHBmslave10_HADDR(19) => 
        CoreAHBLite_0_AHBmslave10_HADDR(19), 
        CoreAHBLite_0_AHBmslave10_HADDR(18) => 
        CoreAHBLite_0_AHBmslave10_HADDR(18), 
        CoreAHBLite_0_AHBmslave10_HADDR(17) => 
        CoreAHBLite_0_AHBmslave10_HADDR(17), 
        CoreAHBLite_0_AHBmslave10_HADDR(16) => 
        CoreAHBLite_0_AHBmslave10_HADDR(16), 
        CoreAHBLite_0_AHBmslave10_HADDR(15) => 
        CoreAHBLite_0_AHBmslave10_HADDR(15), 
        CoreAHBLite_0_AHBmslave10_HADDR(14) => 
        CoreAHBLite_0_AHBmslave10_HADDR(14), 
        CoreAHBLite_0_AHBmslave10_HADDR(13) => 
        CoreAHBLite_0_AHBmslave10_HADDR(13), 
        CoreAHBLite_0_AHBmslave10_HADDR(12) => 
        CoreAHBLite_0_AHBmslave10_HADDR(12), 
        CoreAHBLite_0_AHBmslave10_HADDR(11) => 
        CoreAHBLite_0_AHBmslave10_HADDR(11), 
        CoreAHBLite_0_AHBmslave10_HADDR(10) => 
        CoreAHBLite_0_AHBmslave10_HADDR(10), 
        CoreAHBLite_0_AHBmslave10_HADDR(9) => 
        CoreAHBLite_0_AHBmslave10_HADDR(9), 
        CoreAHBLite_0_AHBmslave10_HADDR(8) => 
        CoreAHBLite_0_AHBmslave10_HADDR(8), 
        CoreAHBLite_0_AHBmslave10_HADDR(7) => 
        CoreAHBLite_0_AHBmslave10_HADDR(7), 
        CoreAHBLite_0_AHBmslave10_HADDR(6) => 
        CoreAHBLite_0_AHBmslave10_HADDR(6), 
        CoreAHBLite_0_AHBmslave10_HADDR(5) => 
        CoreAHBLite_0_AHBmslave10_HADDR(5), 
        CoreAHBLite_0_AHBmslave10_HADDR(4) => 
        CoreAHBLite_0_AHBmslave10_HADDR(4), 
        CoreAHBLite_0_AHBmslave10_HADDR(3) => 
        CoreAHBLite_0_AHBmslave10_HADDR(3), 
        CoreAHBLite_0_AHBmslave10_HADDR(2) => 
        CoreAHBLite_0_AHBmslave10_HADDR(2), 
        CoreAHBLite_0_AHBmslave10_HADDR(1) => 
        CoreAHBLite_0_AHBmslave10_HADDR(1), 
        CoreAHBLite_0_AHBmslave10_HADDR(0) => 
        CoreAHBLite_0_AHBmslave10_HADDR(0), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), xhdl1222_0
         => xhdl1222_0, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0 => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, 
        current_state_0 => current_state_0, masterAddrInProg_0
         => masterAddrInProg_0, hsel2_0_a2_1 => hsel2_0_a2_1, 
        hsel2 => hsel2, CoreAHBLite_0_AHBmslave10_HWRITE => 
        CoreAHBLite_0_AHBmslave10_HWRITE, 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK => 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, MSS_READY => 
        MSS_READY, SDRCLK_c => SDRCLK_c, m0PrevDataSlaveReady => 
        m0PrevDataSlaveReady, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        hready_m_xhdl349 => hready_m_xhdl349, N_91 => N_91, N_92
         => N_92, top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top_sb_CCC_0_FCCC is

    port( FAB_CCC_LOCK : out   std_logic;
          CLK1_PAD     : in    std_logic;
          SDRCLK_c     : out   std_logic
        );

end top_sb_CCC_0_FCCC;

architecture DEF_ARCH of top_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL2_net, CLK1_PAD_net, VCC_net_1, GND_net_1
         : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CLK1_PAD_INST : INBUF
      port map(PAD => CLK1_PAD, Y => CLK1_PAD_net);
    
    GL2_INST : CLKINT
      port map(A => GL2_net, Y => SDRCLK_c);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007F98000044D74000318C1F18C6318C61C40404040401802",
         VCOFREQUENCY => 800.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => CLK1_PAD_net, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => OPEN, GL1
         => OPEN, GL2 => GL2_net, GL3 => OPEN, RCOSC_25_50MHZ => 
        GND_net_1, RCOSC_1MHZ => GND_net_1, XTLOSC => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top_sb_MSS is

    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : out   std_logic_vector(1 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HRDATA              : in    std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : in    std_logic;
          SDRCLK_c                                      : in    std_logic;
          CORERESETP_0_RESET_N_F2M                      : in    std_logic;
          FAB_CCC_LOCK                                  : in    std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : out   std_logic;
          top_sb_MSS_TMP_0_MSS_RESET_N_M2F              : out   std_logic;
          top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N         : out   std_logic;
          hready_m_xhdl349                              : in    std_logic;
          CAN_RX                                        : in    std_logic;
          CAN_TX_EN_N                                   : out   std_logic;
          CAN_TX                                        : out   std_logic;
          GPIO_1_BI                                     : inout std_logic := 'Z';
          GPIO_8_BI                                     : inout std_logic := 'Z';
          GPIO_9_BI                                     : inout std_logic := 'Z';
          GPIO_10_BI                                    : inout std_logic := 'Z';
          GPIO_11_BI                                    : inout std_logic := 'Z';
          GPIO_12_BI                                    : inout std_logic := 'Z';
          GPIO_13_BI                                    : inout std_logic := 'Z';
          GPIO_14_BI                                    : inout std_logic := 'Z';
          GPIO_15_BI                                    : inout std_logic := 'Z';
          GPIO_16_BI                                    : inout std_logic := 'Z';
          GPIO_17_BI                                    : inout std_logic := 'Z';
          GPIO_18_BI                                    : inout std_logic := 'Z';
          GPIO_19_BI                                    : inout std_logic := 'Z';
          GPIO_20_BI                                    : inout std_logic := 'Z';
          GPIO_21_BI                                    : inout std_logic := 'Z';
          GPIO_22_BI                                    : inout std_logic := 'Z';
          GPIO_23_BI                                    : inout std_logic := 'Z';
          GPIO_24_BI                                    : inout std_logic := 'Z';
          GPIO_25_BI                                    : inout std_logic := 'Z';
          GPIO_26_BI                                    : inout std_logic := 'Z';
          GPIO_29_BI                                    : inout std_logic := 'Z';
          I2C_0_SCL                                     : inout std_logic := 'Z';
          I2C_0_SDA                                     : inout std_logic := 'Z';
          MMUART_0_RXD                                  : in    std_logic;
          MMUART_0_TXD                                  : out   std_logic;
          SPI_0_CLK                                     : inout std_logic := 'Z';
          SPI_0_DI                                      : in    std_logic;
          SPI_0_DO                                      : out   std_logic;
          SPI_0_SS0                                     : inout std_logic := 'Z'
        );

end top_sb_MSS;

architecture DEF_ARCH of top_sb_MSS is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component MSS_010

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic
        );
  end component;

    signal SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, I2C_0_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C_0_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE, 
        GPIO_GPIO_29_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OE, 
        GPIO_GPIO_26_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, 
        GPIO_GPIO_25_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, 
        GPIO_GPIO_24_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OUT, 
        MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OE, 
        GPIO_GPIO_23_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OUT, 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OE, 
        GPIO_GPIO_22_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OUT, 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OE, 
        GPIO_GPIO_21_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OUT, 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OE, 
        GPIO_GPIO_20_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OUT, 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OE, 
        GPIO_GPIO_19_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, 
        GPIO_GPIO_18_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        GPIO_GPIO_17_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, 
        GPIO_GPIO_16_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OUT, 
        MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OE, 
        GPIO_GPIO_15_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OUT, 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OE, 
        GPIO_GPIO_14_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OUT, 
        MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OE, 
        GPIO_GPIO_13_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT, 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE, 
        GPIO_GPIO_12_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE, 
        GPIO_GPIO_11_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OUT, 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OE, 
        GPIO_GPIO_10_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OE, 
        GPIO_GPIO_9_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OE, 
        GPIO_GPIO_8_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        GPIO_GPIO_1_BI_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_RX_PAD_Y, \CoreAHBLite_0_AHBmslave10_HRDATA_m[31]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[30]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[29]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[28]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[27]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[26]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[25]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[24]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[23]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[22]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[21]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[20]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[19]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[18]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[17]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[16]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[15]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[14]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[13]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[12]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[11]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[10]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[9]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[8]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[7]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[6]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[5]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[4]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[3]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[2]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[1]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[0]\, VCC_net_1, 
        GND_net_1 : std_logic;
    signal nc228, nc203, nc265, nc216, nc194, nc151, nc23, nc175, 
        nc250, nc58, nc116, nc74, nc133, nc238, nc167, nc84, nc39, 
        nc72, nc256, nc212, nc205, nc82, nc145, nc181, nc160, 
        nc57, nc156, nc280, nc125, nc211, nc73, nc107, nc66, nc83, 
        nc9, nc252, nc171, nc54, nc286, nc307, nc135, nc41, nc100, 
        nc270, nc52, nc251, nc186, nc29, nc269, nc118, nc60, 
        nc141, nc276, nc193, nc214, nc298, nc282, nc240, nc45, 
        nc53, nc121, nc176, nc220, nc158, nc281, nc209, nc246, 
        nc162, nc11, nc272, nc131, nc254, nc267, nc96, nc79, 
        nc226, nc146, nc230, nc89, nc119, nc48, nc271, nc213, 
        nc300, nc126, nc195, nc188, nc242, nc15, nc308, nc236, 
        nc102, nc304, nc3, nc207, nc47, nc90, nc284, nc222, nc159, 
        nc136, nc241, nc253, nc178, nc306, nc215, nc59, nc221, 
        nc232, nc274, nc18, nc44, nc117, nc189, nc164, nc148, 
        nc42, nc231, nc191, nc255, nc283, nc290, nc17, nc2, nc302, 
        nc110, nc128, nc244, nc43, nc179, nc157, nc36, nc224, 
        nc296, nc273, nc61, nc104, nc138, nc14, nc285, nc303, 
        nc150, nc196, nc234, nc149, nc12, nc219, nc30, nc243, 
        nc187, nc65, nc7, nc292, nc129, nc275, nc8, nc223, nc13, 
        nc305, nc180, nc26, nc291, nc177, nc139, nc259, nc245, 
        nc233, nc163, nc268, nc112, nc68, nc49, nc217, nc170, 
        nc91, nc225, nc5, nc20, nc198, nc147, nc67, nc289, nc294, 
        nc152, nc127, nc103, nc235, nc76, nc208, nc140, nc257, 
        nc86, nc95, nc120, nc165, nc279, nc137, nc64, nc19, nc70, 
        nc182, nc62, nc199, nc80, nc130, nc287, nc98, nc293, 
        nc249, nc114, nc56, nc105, nc63, nc172, nc229, nc277, 
        nc97, nc161, nc31, nc295, nc154, nc50, nc260, nc239, 
        nc142, nc247, nc94, nc197, nc122, nc266, nc35, nc4, nc227, 
        nc92, nc101, nc184, nc200, nc190, nc166, nc132, nc21, 
        nc237, nc93, nc262, nc69, nc206, nc174, nc38, nc113, 
        nc218, nc106, nc261, nc25, nc1, nc299, nc37, nc202, nc144, 
        nc153, nc46, nc258, nc71, nc124, nc81, nc201, nc168, nc34, 
        nc28, nc115, nc264, nc192, nc134, nc32, nc40, nc297, nc99, 
        nc75, nc183, nc288, nc85, nc27, nc108, nc16, nc155, nc51, 
        nc301, nc33, nc204, nc173, nc278, nc169, nc78, nc263, 
        nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, 
        nc248, nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 


    MMUART_0_RXD_PAD : INBUF
      port map(PAD => MMUART_0_RXD, Y => MMUART_0_RXD_PAD_Y);
    
    MSS_ADLIB_INST_RNO_20 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(21), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[21]\);
    
    GPIO_GPIO_13_BI_PAD : BIBUF
      port map(PAD => GPIO_13_BI, D => 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE, Y => 
        GPIO_GPIO_13_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_23 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(24), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[24]\);
    
    MSS_ADLIB_INST_RNO_29 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(30), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[30]\);
    
    MSS_ADLIB_INST_RNO_21 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(22), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[22]\);
    
    GPIO_GPIO_25_BI_PAD : BIBUF
      port map(PAD => GPIO_25_BI, D => 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, Y => 
        GPIO_GPIO_25_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(0), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[0]\);
    
    MSS_ADLIB_INST_RNO_22 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(23), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[23]\);
    
    GPIO_GPIO_17_BI_PAD : BIBUF
      port map(PAD => GPIO_17_BI, D => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, Y => 
        GPIO_GPIO_17_BI_PAD_Y);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    GPIO_GPIO_11_BI_PAD : BIBUF
      port map(PAD => GPIO_11_BI, D => 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OE, Y => 
        GPIO_GPIO_11_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_27 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(28), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[28]\);
    
    MSS_ADLIB_INST_RNO_10 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(11), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[11]\);
    
    MMUART_0_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, PAD => 
        MMUART_0_TXD);
    
    GPIO_GPIO_9_BI_PAD : BIBUF
      port map(PAD => GPIO_9_BI, D => 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OE, Y => 
        GPIO_GPIO_9_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_13 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(14), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[14]\);
    
    MSS_ADLIB_INST_RNO_19 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(20), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[20]\);
    
    GPIO_GPIO_23_BI_PAD : BIBUF
      port map(PAD => GPIO_23_BI, D => 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OE, Y => 
        GPIO_GPIO_23_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_11 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(12), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[12]\);
    
    GPIO_GPIO_12_BI_PAD : BIBUF
      port map(PAD => GPIO_12_BI, D => 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE, Y => 
        GPIO_GPIO_12_BI_PAD_Y);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    MSS_ADLIB_INST_RNO_12 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(13), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[13]\);
    
    MSS_ADLIB_INST_RNO_2 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(3), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[3]\);
    
    I2C_0_SCL_PAD : BIBUF
      port map(PAD => I2C_0_SCL, D => 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, E => 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE, Y => 
        I2C_0_SCL_PAD_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    MSS_ADLIB_INST_RNO_4 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(5), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[5]\);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_17 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(18), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[18]\);
    
    CAN_TX_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, E => 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, PAD => 
        CAN_TX);
    
    GPIO_GPIO_21_BI_PAD : BIBUF
      port map(PAD => GPIO_21_BI, D => 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OE, Y => 
        GPIO_GPIO_21_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_7 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(8), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[8]\);
    
    GPIO_GPIO_1_BI_PAD : BIBUF
      port map(PAD => GPIO_1_BI, D => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, Y => 
        GPIO_GPIO_1_BI_PAD_Y);
    
    GPIO_GPIO_14_BI_PAD : BIBUF
      port map(PAD => GPIO_14_BI, D => 
        MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OE, Y => 
        GPIO_GPIO_14_BI_PAD_Y);
    
    MSS_ADLIB_INST : MSS_010

              generic map(INIT => "00" & x"000040190B612024290A4290800002429080000000000000000090A4290A4290A4290A4290A42000000000090A4290801203612036120242000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000200006092C0104003FFFFE0000000000020326780000F0F01C000000025544010842108421000001FE34001FF8000000480000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 100.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => OPEN, COMMS_INT => OPEN, 
        CONFIG_PRESET_N => top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc265, EDAC_ERROR(4) => nc216, 
        EDAC_ERROR(3) => nc194, EDAC_ERROR(2) => nc151, 
        EDAC_ERROR(1) => nc23, EDAC_ERROR(0) => nc175, 
        F_FM0_RDATA(31) => nc250, F_FM0_RDATA(30) => nc58, 
        F_FM0_RDATA(29) => nc116, F_FM0_RDATA(28) => nc74, 
        F_FM0_RDATA(27) => nc133, F_FM0_RDATA(26) => nc238, 
        F_FM0_RDATA(25) => nc167, F_FM0_RDATA(24) => nc84, 
        F_FM0_RDATA(23) => nc39, F_FM0_RDATA(22) => nc72, 
        F_FM0_RDATA(21) => nc256, F_FM0_RDATA(20) => nc212, 
        F_FM0_RDATA(19) => nc205, F_FM0_RDATA(18) => nc82, 
        F_FM0_RDATA(17) => nc145, F_FM0_RDATA(16) => nc181, 
        F_FM0_RDATA(15) => nc160, F_FM0_RDATA(14) => nc57, 
        F_FM0_RDATA(13) => nc156, F_FM0_RDATA(12) => nc280, 
        F_FM0_RDATA(11) => nc125, F_FM0_RDATA(10) => nc211, 
        F_FM0_RDATA(9) => nc73, F_FM0_RDATA(8) => nc107, 
        F_FM0_RDATA(7) => nc66, F_FM0_RDATA(6) => nc83, 
        F_FM0_RDATA(5) => nc9, F_FM0_RDATA(4) => nc252, 
        F_FM0_RDATA(3) => nc171, F_FM0_RDATA(2) => nc54, 
        F_FM0_RDATA(1) => nc286, F_FM0_RDATA(0) => nc307, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc135, F_HM0_ADDR(30) => nc41, 
        F_HM0_ADDR(29) => nc100, F_HM0_ADDR(28) => nc270, 
        F_HM0_ADDR(27) => nc52, F_HM0_ADDR(26) => nc251, 
        F_HM0_ADDR(25) => nc186, F_HM0_ADDR(24) => nc29, 
        F_HM0_ADDR(23) => nc269, F_HM0_ADDR(22) => nc118, 
        F_HM0_ADDR(21) => nc60, F_HM0_ADDR(20) => nc141, 
        F_HM0_ADDR(19) => nc276, F_HM0_ADDR(18) => nc193, 
        F_HM0_ADDR(17) => nc214, F_HM0_ADDR(16) => nc298, 
        F_HM0_ADDR(15) => nc282, F_HM0_ADDR(14) => nc240, 
        F_HM0_ADDR(13) => nc45, F_HM0_ADDR(12) => nc53, 
        F_HM0_ADDR(11) => nc121, F_HM0_ADDR(10) => nc176, 
        F_HM0_ADDR(9) => nc220, F_HM0_ADDR(8) => nc158, 
        F_HM0_ADDR(7) => nc281, F_HM0_ADDR(6) => nc209, 
        F_HM0_ADDR(5) => nc246, F_HM0_ADDR(4) => nc162, 
        F_HM0_ADDR(3) => nc11, F_HM0_ADDR(2) => nc272, 
        F_HM0_ADDR(1) => nc131, F_HM0_ADDR(0) => nc254, 
        F_HM0_ENABLE => OPEN, F_HM0_SEL => OPEN, F_HM0_SIZE(1)
         => nc267, F_HM0_SIZE(0) => nc96, F_HM0_TRANS1 => OPEN, 
        F_HM0_WDATA(31) => nc79, F_HM0_WDATA(30) => nc226, 
        F_HM0_WDATA(29) => nc146, F_HM0_WDATA(28) => nc230, 
        F_HM0_WDATA(27) => nc89, F_HM0_WDATA(26) => nc119, 
        F_HM0_WDATA(25) => nc48, F_HM0_WDATA(24) => nc271, 
        F_HM0_WDATA(23) => nc213, F_HM0_WDATA(22) => nc300, 
        F_HM0_WDATA(21) => nc126, F_HM0_WDATA(20) => nc195, 
        F_HM0_WDATA(19) => nc188, F_HM0_WDATA(18) => nc242, 
        F_HM0_WDATA(17) => nc15, F_HM0_WDATA(16) => nc308, 
        F_HM0_WDATA(15) => nc236, F_HM0_WDATA(14) => nc102, 
        F_HM0_WDATA(13) => nc304, F_HM0_WDATA(12) => nc3, 
        F_HM0_WDATA(11) => nc207, F_HM0_WDATA(10) => nc47, 
        F_HM0_WDATA(9) => nc90, F_HM0_WDATA(8) => nc284, 
        F_HM0_WDATA(7) => nc222, F_HM0_WDATA(6) => nc159, 
        F_HM0_WDATA(5) => nc136, F_HM0_WDATA(4) => nc241, 
        F_HM0_WDATA(3) => nc253, F_HM0_WDATA(2) => nc178, 
        F_HM0_WDATA(1) => nc306, F_HM0_WDATA(0) => nc215, 
        F_HM0_WRITE => OPEN, FAB_CHRGVBUS => OPEN, 
        FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc59, FAB_OPMODE(0) => nc221, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc232, FAB_VCONTROL(2) => 
        nc274, FAB_VCONTROL(1) => nc18, FAB_VCONTROL(0) => nc44, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc117, 
        FAB_XCVRSEL(0) => nc189, FAB_XDATAOUT(7) => nc164, 
        FAB_XDATAOUT(6) => nc148, FAB_XDATAOUT(5) => nc42, 
        FAB_XDATAOUT(4) => nc231, FAB_XDATAOUT(3) => nc191, 
        FAB_XDATAOUT(2) => nc255, FAB_XDATAOUT(1) => nc283, 
        FAB_XDATAOUT(0) => nc290, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc17, FIC32_0_MASTER(0) => nc2, 
        FIC32_1_MASTER(1) => nc302, FIC32_1_MASTER(0) => nc110, 
        FPGA_RESET_N => top_sb_MSS_TMP_0_MSS_RESET_N_M2F, GTX_CLK
         => OPEN, H2F_INTERRUPT(15) => nc128, H2F_INTERRUPT(14)
         => nc244, H2F_INTERRUPT(13) => nc43, H2F_INTERRUPT(12)
         => nc179, H2F_INTERRUPT(11) => nc157, H2F_INTERRUPT(10)
         => nc36, H2F_INTERRUPT(9) => nc224, H2F_INTERRUPT(8) => 
        nc296, H2F_INTERRUPT(7) => nc273, H2F_INTERRUPT(6) => 
        nc61, H2F_INTERRUPT(5) => nc104, H2F_INTERRUPT(4) => 
        nc138, H2F_INTERRUPT(3) => nc14, H2F_INTERRUPT(2) => 
        nc285, H2F_INTERRUPT(1) => nc303, H2F_INTERRUPT(0) => 
        nc150, H2F_NMI => OPEN, H2FCALIB => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_A => OPEN, I2C0_SCL_MGPIO31B_H2F_B
         => OPEN, I2C0_SDA_MGPIO30B_H2F_A => OPEN, 
        I2C0_SDA_MGPIO30B_H2F_B => OPEN, I2C1_SCL_MGPIO1A_H2F_A
         => OPEN, I2C1_SCL_MGPIO1A_H2F_B => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_A => OPEN, I2C1_SDA_MGPIO0A_H2F_B
         => OPEN, MDCF => OPEN, MDOENF => OPEN, MDOF => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => OPEN, MPLL_LOCK => OPEN, 
        PER2_FABRIC_PADDR(15) => nc196, PER2_FABRIC_PADDR(14) => 
        nc234, PER2_FABRIC_PADDR(13) => nc149, 
        PER2_FABRIC_PADDR(12) => nc12, PER2_FABRIC_PADDR(11) => 
        nc219, PER2_FABRIC_PADDR(10) => nc30, 
        PER2_FABRIC_PADDR(9) => nc243, PER2_FABRIC_PADDR(8) => 
        nc187, PER2_FABRIC_PADDR(7) => nc65, PER2_FABRIC_PADDR(6)
         => nc7, PER2_FABRIC_PADDR(5) => nc292, 
        PER2_FABRIC_PADDR(4) => nc129, PER2_FABRIC_PADDR(3) => 
        nc275, PER2_FABRIC_PADDR(2) => nc8, PER2_FABRIC_PENABLE
         => OPEN, PER2_FABRIC_PSEL => OPEN, 
        PER2_FABRIC_PWDATA(31) => nc223, PER2_FABRIC_PWDATA(30)
         => nc13, PER2_FABRIC_PWDATA(29) => nc305, 
        PER2_FABRIC_PWDATA(28) => nc180, PER2_FABRIC_PWDATA(27)
         => nc26, PER2_FABRIC_PWDATA(26) => nc291, 
        PER2_FABRIC_PWDATA(25) => nc177, PER2_FABRIC_PWDATA(24)
         => nc139, PER2_FABRIC_PWDATA(23) => nc259, 
        PER2_FABRIC_PWDATA(22) => nc245, PER2_FABRIC_PWDATA(21)
         => nc233, PER2_FABRIC_PWDATA(20) => nc163, 
        PER2_FABRIC_PWDATA(19) => nc268, PER2_FABRIC_PWDATA(18)
         => nc112, PER2_FABRIC_PWDATA(17) => nc68, 
        PER2_FABRIC_PWDATA(16) => nc49, PER2_FABRIC_PWDATA(15)
         => nc217, PER2_FABRIC_PWDATA(14) => nc170, 
        PER2_FABRIC_PWDATA(13) => nc91, PER2_FABRIC_PWDATA(12)
         => nc225, PER2_FABRIC_PWDATA(11) => nc5, 
        PER2_FABRIC_PWDATA(10) => nc20, PER2_FABRIC_PWDATA(9) => 
        nc198, PER2_FABRIC_PWDATA(8) => nc147, 
        PER2_FABRIC_PWDATA(7) => nc67, PER2_FABRIC_PWDATA(6) => 
        nc289, PER2_FABRIC_PWDATA(5) => nc294, 
        PER2_FABRIC_PWDATA(4) => nc152, PER2_FABRIC_PWDATA(3) => 
        nc127, PER2_FABRIC_PWDATA(2) => nc103, 
        PER2_FABRIC_PWDATA(1) => nc235, PER2_FABRIC_PWDATA(0) => 
        nc76, PER2_FABRIC_PWRITE => OPEN, RTC_MATCH => OPEN, 
        SLEEPDEEP => OPEN, SLEEPHOLDACK => OPEN, SLEEPING => OPEN, 
        SMBALERT_NO0 => OPEN, SMBALERT_NO1 => OPEN, SMBSUS_NO0
         => OPEN, SMBSUS_NO1 => OPEN, SPI0_CLK_OUT => OPEN, 
        SPI0_SDI_MGPIO5A_H2F_A => OPEN, SPI0_SDI_MGPIO5A_H2F_B
         => OPEN, SPI0_SDO_MGPIO6A_H2F_A => OPEN, 
        SPI0_SDO_MGPIO6A_H2F_B => OPEN, SPI0_SS0_MGPIO7A_H2F_A
         => OPEN, SPI0_SS0_MGPIO7A_H2F_B => OPEN, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => OPEN, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => OPEN, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => OPEN, SPI1_SDO_MGPIO12A_H2F_A => OPEN, 
        SPI1_SDO_MGPIO12A_H2F_B => OPEN, SPI1_SS0_MGPIO13A_H2F_A
         => OPEN, SPI1_SS0_MGPIO13A_H2F_B => OPEN, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc208, 
        TCGF(8) => nc140, TCGF(7) => nc257, TCGF(6) => nc86, 
        TCGF(5) => nc95, TCGF(4) => nc120, TCGF(3) => nc165, 
        TCGF(2) => nc279, TCGF(1) => nc137, TCGF(0) => nc64, 
        TRACECLK => OPEN, TRACEDATA(3) => nc19, TRACEDATA(2) => 
        nc70, TRACEDATA(1) => nc182, TRACEDATA(0) => nc62, TX_CLK
         => OPEN, TX_ENF => OPEN, TX_ERRF => OPEN, TXCTL_EN_RIF
         => OPEN, TXD_RIF(3) => nc199, TXD_RIF(2) => nc80, 
        TXD_RIF(1) => nc130, TXD_RIF(0) => nc287, TXDF(7) => nc98, 
        TXDF(6) => nc293, TXDF(5) => nc249, TXDF(4) => nc114, 
        TXDF(3) => nc56, TXDF(2) => nc105, TXDF(1) => nc63, 
        TXDF(0) => nc172, TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        F_AWREADY_HREADYOUT0 => OPEN, F_BID(3) => nc229, F_BID(2)
         => nc277, F_BID(1) => nc97, F_BID(0) => nc161, 
        F_BRESP_HRESP0(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0, 
        F_BRESP_HRESP0(0) => nc31, F_BVALID => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        F_RDATA_HRDATA01(63) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31), 
        F_RDATA_HRDATA01(62) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30), 
        F_RDATA_HRDATA01(61) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29), 
        F_RDATA_HRDATA01(60) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28), 
        F_RDATA_HRDATA01(59) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27), 
        F_RDATA_HRDATA01(58) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26), 
        F_RDATA_HRDATA01(57) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25), 
        F_RDATA_HRDATA01(56) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24), 
        F_RDATA_HRDATA01(55) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23), 
        F_RDATA_HRDATA01(54) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22), 
        F_RDATA_HRDATA01(53) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21), 
        F_RDATA_HRDATA01(52) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20), 
        F_RDATA_HRDATA01(51) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19), 
        F_RDATA_HRDATA01(50) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18), 
        F_RDATA_HRDATA01(49) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17), 
        F_RDATA_HRDATA01(48) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16), 
        F_RDATA_HRDATA01(47) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15), 
        F_RDATA_HRDATA01(46) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14), 
        F_RDATA_HRDATA01(45) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13), 
        F_RDATA_HRDATA01(44) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12), 
        F_RDATA_HRDATA01(43) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11), 
        F_RDATA_HRDATA01(42) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10), 
        F_RDATA_HRDATA01(41) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9), 
        F_RDATA_HRDATA01(40) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8), 
        F_RDATA_HRDATA01(39) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7), 
        F_RDATA_HRDATA01(38) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6), 
        F_RDATA_HRDATA01(37) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5), 
        F_RDATA_HRDATA01(36) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4), 
        F_RDATA_HRDATA01(35) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3), 
        F_RDATA_HRDATA01(34) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2), 
        F_RDATA_HRDATA01(33) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1), 
        F_RDATA_HRDATA01(32) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0), 
        F_RDATA_HRDATA01(31) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31), 
        F_RDATA_HRDATA01(30) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30), 
        F_RDATA_HRDATA01(29) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29), 
        F_RDATA_HRDATA01(28) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28), 
        F_RDATA_HRDATA01(27) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27), 
        F_RDATA_HRDATA01(26) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26), 
        F_RDATA_HRDATA01(25) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25), 
        F_RDATA_HRDATA01(24) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24), 
        F_RDATA_HRDATA01(23) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23), 
        F_RDATA_HRDATA01(22) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22), 
        F_RDATA_HRDATA01(21) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21), 
        F_RDATA_HRDATA01(20) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20), 
        F_RDATA_HRDATA01(19) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19), 
        F_RDATA_HRDATA01(18) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18), 
        F_RDATA_HRDATA01(17) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17), 
        F_RDATA_HRDATA01(16) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16), 
        F_RDATA_HRDATA01(15) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15), 
        F_RDATA_HRDATA01(14) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14), 
        F_RDATA_HRDATA01(13) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13), 
        F_RDATA_HRDATA01(12) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12), 
        F_RDATA_HRDATA01(11) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11), 
        F_RDATA_HRDATA01(10) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10), 
        F_RDATA_HRDATA01(9) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9), 
        F_RDATA_HRDATA01(8) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8), 
        F_RDATA_HRDATA01(7) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7), 
        F_RDATA_HRDATA01(6) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6), 
        F_RDATA_HRDATA01(5) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5), 
        F_RDATA_HRDATA01(4) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4), 
        F_RDATA_HRDATA01(3) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3), 
        F_RDATA_HRDATA01(2) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2), 
        F_RDATA_HRDATA01(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1), 
        F_RDATA_HRDATA01(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0), F_RID(3)
         => nc295, F_RID(2) => nc154, F_RID(1) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1), F_RID(0)
         => top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0), 
        F_RLAST => OPEN, F_RRESP_HRESP1(1) => nc50, 
        F_RRESP_HRESP1(0) => nc260, F_RVALID => OPEN, F_WREADY
         => OPEN, MDDR_FABRIC_PRDATA(15) => nc239, 
        MDDR_FABRIC_PRDATA(14) => nc142, MDDR_FABRIC_PRDATA(13)
         => nc247, MDDR_FABRIC_PRDATA(12) => nc94, 
        MDDR_FABRIC_PRDATA(11) => nc197, MDDR_FABRIC_PRDATA(10)
         => nc122, MDDR_FABRIC_PRDATA(9) => nc266, 
        MDDR_FABRIC_PRDATA(8) => nc35, MDDR_FABRIC_PRDATA(7) => 
        nc4, MDDR_FABRIC_PRDATA(6) => nc227, 
        MDDR_FABRIC_PRDATA(5) => nc92, MDDR_FABRIC_PRDATA(4) => 
        nc101, MDDR_FABRIC_PRDATA(3) => nc184, 
        MDDR_FABRIC_PRDATA(2) => nc200, MDDR_FABRIC_PRDATA(1) => 
        nc190, MDDR_FABRIC_PRDATA(0) => nc166, MDDR_FABRIC_PREADY
         => OPEN, MDDR_FABRIC_PSLVERR => OPEN, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => VCC_net_1, CRSF
         => VCC_net_1, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        GND_net_1, F2HCALIB => VCC_net_1, F_DMAREADY(1) => 
        VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31) => 
        GND_net_1, F_FM0_ADDR(30) => GND_net_1, F_FM0_ADDR(29)
         => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => GND_net_1, F_HM0_RDATA(30) => 
        GND_net_1, F_HM0_RDATA(29) => GND_net_1, F_HM0_RDATA(28)
         => GND_net_1, F_HM0_RDATA(27) => GND_net_1, 
        F_HM0_RDATA(26) => GND_net_1, F_HM0_RDATA(25) => 
        GND_net_1, F_HM0_RDATA(24) => GND_net_1, F_HM0_RDATA(23)
         => GND_net_1, F_HM0_RDATA(22) => GND_net_1, 
        F_HM0_RDATA(21) => GND_net_1, F_HM0_RDATA(20) => 
        GND_net_1, F_HM0_RDATA(19) => GND_net_1, F_HM0_RDATA(18)
         => GND_net_1, F_HM0_RDATA(17) => GND_net_1, 
        F_HM0_RDATA(16) => GND_net_1, F_HM0_RDATA(15) => 
        GND_net_1, F_HM0_RDATA(14) => GND_net_1, F_HM0_RDATA(13)
         => GND_net_1, F_HM0_RDATA(12) => GND_net_1, 
        F_HM0_RDATA(11) => GND_net_1, F_HM0_RDATA(10) => 
        GND_net_1, F_HM0_RDATA(9) => GND_net_1, F_HM0_RDATA(8)
         => GND_net_1, F_HM0_RDATA(7) => GND_net_1, 
        F_HM0_RDATA(6) => GND_net_1, F_HM0_RDATA(5) => GND_net_1, 
        F_HM0_RDATA(4) => GND_net_1, F_HM0_RDATA(3) => GND_net_1, 
        F_HM0_RDATA(2) => GND_net_1, F_HM0_RDATA(1) => GND_net_1, 
        F_HM0_RDATA(0) => GND_net_1, F_HM0_READY => VCC_net_1, 
        F_HM0_RESP => GND_net_1, FAB_AVALID => VCC_net_1, 
        FAB_HOSTDISCON => VCC_net_1, FAB_IDDIG => VCC_net_1, 
        FAB_LINESTATE(1) => VCC_net_1, FAB_LINESTATE(0) => 
        VCC_net_1, FAB_M3_RESET_N => VCC_net_1, FAB_PLL_LOCK => 
        FAB_CCC_LOCK, FAB_RXACTIVE => VCC_net_1, FAB_RXERROR => 
        VCC_net_1, FAB_RXVALID => VCC_net_1, FAB_RXVALIDH => 
        GND_net_1, FAB_SESSEND => VCC_net_1, FAB_TXREADY => 
        VCC_net_1, FAB_VBUSVALID => VCC_net_1, FAB_VSTATUS(7) => 
        VCC_net_1, FAB_VSTATUS(6) => VCC_net_1, FAB_VSTATUS(5)
         => VCC_net_1, FAB_VSTATUS(4) => VCC_net_1, 
        FAB_VSTATUS(3) => VCC_net_1, FAB_VSTATUS(2) => VCC_net_1, 
        FAB_VSTATUS(1) => VCC_net_1, FAB_VSTATUS(0) => VCC_net_1, 
        FAB_XDATAIN(7) => VCC_net_1, FAB_XDATAIN(6) => VCC_net_1, 
        FAB_XDATAIN(5) => VCC_net_1, FAB_XDATAIN(4) => VCC_net_1, 
        FAB_XDATAIN(3) => VCC_net_1, FAB_XDATAIN(2) => VCC_net_1, 
        FAB_XDATAIN(1) => VCC_net_1, FAB_XDATAIN(0) => VCC_net_1, 
        GTX_CLKPF => VCC_net_1, I2C0_BCLK => VCC_net_1, 
        I2C0_SCL_F2H_SCP => VCC_net_1, I2C0_SDA_F2H_SCP => 
        VCC_net_1, I2C1_BCLK => VCC_net_1, I2C1_SCL_F2H_SCP => 
        VCC_net_1, I2C1_SDA_F2H_SCP => VCC_net_1, MDIF => 
        VCC_net_1, MGPIO0A_F2H_GPIN => VCC_net_1, 
        MGPIO10A_F2H_GPIN => VCC_net_1, MGPIO11A_F2H_GPIN => 
        VCC_net_1, MGPIO11B_F2H_GPIN => VCC_net_1, 
        MGPIO12A_F2H_GPIN => VCC_net_1, MGPIO13A_F2H_GPIN => 
        VCC_net_1, MGPIO14A_F2H_GPIN => VCC_net_1, 
        MGPIO15A_F2H_GPIN => VCC_net_1, MGPIO16A_F2H_GPIN => 
        VCC_net_1, MGPIO17B_F2H_GPIN => VCC_net_1, 
        MGPIO18B_F2H_GPIN => VCC_net_1, MGPIO19B_F2H_GPIN => 
        VCC_net_1, MGPIO1A_F2H_GPIN => VCC_net_1, 
        MGPIO20B_F2H_GPIN => VCC_net_1, MGPIO21B_F2H_GPIN => 
        VCC_net_1, MGPIO22B_F2H_GPIN => VCC_net_1, 
        MGPIO24B_F2H_GPIN => VCC_net_1, MGPIO25B_F2H_GPIN => 
        VCC_net_1, MGPIO26B_F2H_GPIN => VCC_net_1, 
        MGPIO27B_F2H_GPIN => VCC_net_1, MGPIO28B_F2H_GPIN => 
        VCC_net_1, MGPIO29B_F2H_GPIN => VCC_net_1, 
        MGPIO2A_F2H_GPIN => VCC_net_1, MGPIO30B_F2H_GPIN => 
        VCC_net_1, MGPIO31B_F2H_GPIN => VCC_net_1, 
        MGPIO3A_F2H_GPIN => VCC_net_1, MGPIO4A_F2H_GPIN => 
        VCC_net_1, MGPIO5A_F2H_GPIN => VCC_net_1, 
        MGPIO6A_F2H_GPIN => VCC_net_1, MGPIO7A_F2H_GPIN => 
        VCC_net_1, MGPIO8A_F2H_GPIN => VCC_net_1, 
        MGPIO9A_F2H_GPIN => VCC_net_1, MMUART0_CTS_F2H_SCP => 
        VCC_net_1, MMUART0_DCD_F2H_SCP => VCC_net_1, 
        MMUART0_DSR_F2H_SCP => VCC_net_1, MMUART0_DTR_F2H_SCP => 
        VCC_net_1, MMUART0_RI_F2H_SCP => VCC_net_1, 
        MMUART0_RTS_F2H_SCP => VCC_net_1, MMUART0_RXD_F2H_SCP => 
        VCC_net_1, MMUART0_SCK_F2H_SCP => VCC_net_1, 
        MMUART0_TXD_F2H_SCP => VCC_net_1, MMUART1_CTS_F2H_SCP => 
        VCC_net_1, MMUART1_DCD_F2H_SCP => VCC_net_1, 
        MMUART1_DSR_F2H_SCP => VCC_net_1, MMUART1_RI_F2H_SCP => 
        VCC_net_1, MMUART1_RTS_F2H_SCP => VCC_net_1, 
        MMUART1_RXD_F2H_SCP => VCC_net_1, MMUART1_SCK_F2H_SCP => 
        VCC_net_1, MMUART1_TXD_F2H_SCP => VCC_net_1, 
        PER2_FABRIC_PRDATA(31) => GND_net_1, 
        PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => GND_net_1, 
        PER2_FABRIC_PRDATA(17) => GND_net_1, 
        PER2_FABRIC_PRDATA(16) => GND_net_1, 
        PER2_FABRIC_PRDATA(15) => GND_net_1, 
        PER2_FABRIC_PRDATA(14) => GND_net_1, 
        PER2_FABRIC_PRDATA(13) => GND_net_1, 
        PER2_FABRIC_PRDATA(12) => GND_net_1, 
        PER2_FABRIC_PRDATA(11) => GND_net_1, 
        PER2_FABRIC_PRDATA(10) => GND_net_1, 
        PER2_FABRIC_PRDATA(9) => GND_net_1, PER2_FABRIC_PRDATA(8)
         => GND_net_1, PER2_FABRIC_PRDATA(7) => GND_net_1, 
        PER2_FABRIC_PRDATA(6) => GND_net_1, PER2_FABRIC_PRDATA(5)
         => GND_net_1, PER2_FABRIC_PRDATA(4) => GND_net_1, 
        PER2_FABRIC_PRDATA(3) => GND_net_1, PER2_FABRIC_PRDATA(2)
         => GND_net_1, PER2_FABRIC_PRDATA(1) => GND_net_1, 
        PER2_FABRIC_PRDATA(0) => GND_net_1, PER2_FABRIC_PREADY
         => VCC_net_1, PER2_FABRIC_PSLVERR => GND_net_1, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        VCC_net_1, RX_DVF => VCC_net_1, RX_ERRF => VCC_net_1, 
        RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, RXDF(6) => 
        VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => VCC_net_1, 
        RXDF(3) => VCC_net_1, RXDF(2) => VCC_net_1, RXDF(1) => 
        VCC_net_1, RXDF(0) => VCC_net_1, SLEEPHOLDREQ => 
        GND_net_1, SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => 
        VCC_net_1, SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => 
        VCC_net_1, SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => 
        VCC_net_1, SPI0_SDO_F2H_SCP => VCC_net_1, 
        SPI0_SS0_F2H_SCP => VCC_net_1, SPI0_SS1_F2H_SCP => 
        VCC_net_1, SPI0_SS2_F2H_SCP => VCC_net_1, 
        SPI0_SS3_F2H_SCP => VCC_net_1, SPI1_CLK_IN => VCC_net_1, 
        SPI1_SDI_F2H_SCP => VCC_net_1, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => VCC_net_1, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        VCC_net_1, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => CORERESETP_0_RESET_N_F2M, XCLK_FAB
         => VCC_net_1, CLK_BASE => SDRCLK_c, CLK_MDDR_APB => 
        VCC_net_1, F_ARADDR_HADDR1(31) => VCC_net_1, 
        F_ARADDR_HADDR1(30) => VCC_net_1, F_ARADDR_HADDR1(29) => 
        VCC_net_1, F_ARADDR_HADDR1(28) => VCC_net_1, 
        F_ARADDR_HADDR1(27) => VCC_net_1, F_ARADDR_HADDR1(26) => 
        VCC_net_1, F_ARADDR_HADDR1(25) => VCC_net_1, 
        F_ARADDR_HADDR1(24) => VCC_net_1, F_ARADDR_HADDR1(23) => 
        VCC_net_1, F_ARADDR_HADDR1(22) => VCC_net_1, 
        F_ARADDR_HADDR1(21) => VCC_net_1, F_ARADDR_HADDR1(20) => 
        VCC_net_1, F_ARADDR_HADDR1(19) => VCC_net_1, 
        F_ARADDR_HADDR1(18) => VCC_net_1, F_ARADDR_HADDR1(17) => 
        VCC_net_1, F_ARADDR_HADDR1(16) => VCC_net_1, 
        F_ARADDR_HADDR1(15) => VCC_net_1, F_ARADDR_HADDR1(14) => 
        VCC_net_1, F_ARADDR_HADDR1(13) => VCC_net_1, 
        F_ARADDR_HADDR1(12) => VCC_net_1, F_ARADDR_HADDR1(11) => 
        VCC_net_1, F_ARADDR_HADDR1(10) => VCC_net_1, 
        F_ARADDR_HADDR1(9) => VCC_net_1, F_ARADDR_HADDR1(8) => 
        VCC_net_1, F_ARADDR_HADDR1(7) => VCC_net_1, 
        F_ARADDR_HADDR1(6) => VCC_net_1, F_ARADDR_HADDR1(5) => 
        VCC_net_1, F_ARADDR_HADDR1(4) => VCC_net_1, 
        F_ARADDR_HADDR1(3) => VCC_net_1, F_ARADDR_HADDR1(2) => 
        VCC_net_1, F_ARADDR_HADDR1(1) => VCC_net_1, 
        F_ARADDR_HADDR1(0) => VCC_net_1, F_ARBURST_HTRANS1(1) => 
        GND_net_1, F_ARBURST_HTRANS1(0) => GND_net_1, 
        F_ARID_HSEL1(3) => GND_net_1, F_ARID_HSEL1(2) => 
        GND_net_1, F_ARID_HSEL1(1) => GND_net_1, F_ARID_HSEL1(0)
         => GND_net_1, F_ARLEN_HBURST1(3) => GND_net_1, 
        F_ARLEN_HBURST1(2) => GND_net_1, F_ARLEN_HBURST1(1) => 
        GND_net_1, F_ARLEN_HBURST1(0) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(1) => GND_net_1, 
        F_ARLOCK_HMASTLOCK1(0) => GND_net_1, F_ARSIZE_HSIZE1(1)
         => GND_net_1, F_ARSIZE_HSIZE1(0) => GND_net_1, 
        F_ARVALID_HWRITE1 => GND_net_1, F_AWADDR_HADDR0(31) => 
        VCC_net_1, F_AWADDR_HADDR0(30) => VCC_net_1, 
        F_AWADDR_HADDR0(29) => VCC_net_1, F_AWADDR_HADDR0(28) => 
        VCC_net_1, F_AWADDR_HADDR0(27) => VCC_net_1, 
        F_AWADDR_HADDR0(26) => VCC_net_1, F_AWADDR_HADDR0(25) => 
        VCC_net_1, F_AWADDR_HADDR0(24) => VCC_net_1, 
        F_AWADDR_HADDR0(23) => VCC_net_1, F_AWADDR_HADDR0(22) => 
        VCC_net_1, F_AWADDR_HADDR0(21) => VCC_net_1, 
        F_AWADDR_HADDR0(20) => VCC_net_1, F_AWADDR_HADDR0(19) => 
        VCC_net_1, F_AWADDR_HADDR0(18) => VCC_net_1, 
        F_AWADDR_HADDR0(17) => VCC_net_1, F_AWADDR_HADDR0(16) => 
        VCC_net_1, F_AWADDR_HADDR0(15) => VCC_net_1, 
        F_AWADDR_HADDR0(14) => VCC_net_1, F_AWADDR_HADDR0(13) => 
        VCC_net_1, F_AWADDR_HADDR0(12) => VCC_net_1, 
        F_AWADDR_HADDR0(11) => VCC_net_1, F_AWADDR_HADDR0(10) => 
        VCC_net_1, F_AWADDR_HADDR0(9) => VCC_net_1, 
        F_AWADDR_HADDR0(8) => VCC_net_1, F_AWADDR_HADDR0(7) => 
        VCC_net_1, F_AWADDR_HADDR0(6) => VCC_net_1, 
        F_AWADDR_HADDR0(5) => VCC_net_1, F_AWADDR_HADDR0(4) => 
        VCC_net_1, F_AWADDR_HADDR0(3) => VCC_net_1, 
        F_AWADDR_HADDR0(2) => VCC_net_1, F_AWADDR_HADDR0(1) => 
        VCC_net_1, F_AWADDR_HADDR0(0) => VCC_net_1, 
        F_AWBURST_HTRANS0(1) => GND_net_1, F_AWBURST_HTRANS0(0)
         => GND_net_1, F_AWID_HSEL0(3) => GND_net_1, 
        F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1) => 
        GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[31]\, 
        F_WDATA_HWDATA01(30) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[30]\, 
        F_WDATA_HWDATA01(29) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[29]\, 
        F_WDATA_HWDATA01(28) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[28]\, 
        F_WDATA_HWDATA01(27) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[27]\, 
        F_WDATA_HWDATA01(26) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[26]\, 
        F_WDATA_HWDATA01(25) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[25]\, 
        F_WDATA_HWDATA01(24) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[24]\, 
        F_WDATA_HWDATA01(23) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[23]\, 
        F_WDATA_HWDATA01(22) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[22]\, 
        F_WDATA_HWDATA01(21) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[21]\, 
        F_WDATA_HWDATA01(20) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[20]\, 
        F_WDATA_HWDATA01(19) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[19]\, 
        F_WDATA_HWDATA01(18) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[18]\, 
        F_WDATA_HWDATA01(17) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[17]\, 
        F_WDATA_HWDATA01(16) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[16]\, 
        F_WDATA_HWDATA01(15) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[15]\, 
        F_WDATA_HWDATA01(14) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[14]\, 
        F_WDATA_HWDATA01(13) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[13]\, 
        F_WDATA_HWDATA01(12) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[12]\, 
        F_WDATA_HWDATA01(11) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[11]\, 
        F_WDATA_HWDATA01(10) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[10]\, 
        F_WDATA_HWDATA01(9) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[9]\, 
        F_WDATA_HWDATA01(8) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[8]\, 
        F_WDATA_HWDATA01(7) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[7]\, 
        F_WDATA_HWDATA01(6) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[6]\, 
        F_WDATA_HWDATA01(5) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[5]\, 
        F_WDATA_HWDATA01(4) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[4]\, 
        F_WDATA_HWDATA01(3) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[3]\, 
        F_WDATA_HWDATA01(2) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[2]\, 
        F_WDATA_HWDATA01(1) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[1]\, 
        F_WDATA_HWDATA01(0) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[0]\, 
        F_WID_HREADY01(3) => GND_net_1, F_WID_HREADY01(2) => 
        GND_net_1, F_WID_HREADY01(1) => GND_net_1, 
        F_WID_HREADY01(0) => GND_net_1, F_WLAST => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY, F_WSTRB(7)
         => GND_net_1, F_WSTRB(6) => GND_net_1, F_WSTRB(5) => 
        GND_net_1, F_WSTRB(4) => GND_net_1, F_WSTRB(3) => 
        GND_net_1, F_WSTRB(2) => GND_net_1, F_WSTRB(1) => 
        GND_net_1, F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => VCC_net_1, MDDR_FABRIC_PADDR(9) => VCC_net_1, 
        MDDR_FABRIC_PADDR(8) => VCC_net_1, MDDR_FABRIC_PADDR(7)
         => VCC_net_1, MDDR_FABRIC_PADDR(6) => VCC_net_1, 
        MDDR_FABRIC_PADDR(5) => VCC_net_1, MDDR_FABRIC_PADDR(4)
         => VCC_net_1, MDDR_FABRIC_PADDR(3) => VCC_net_1, 
        MDDR_FABRIC_PADDR(2) => VCC_net_1, MDDR_FABRIC_PENABLE
         => VCC_net_1, MDDR_FABRIC_PSEL => VCC_net_1, 
        MDDR_FABRIC_PWDATA(15) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(14) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(13) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(12) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(11) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(10) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(9) => VCC_net_1, MDDR_FABRIC_PWDATA(8)
         => VCC_net_1, MDDR_FABRIC_PWDATA(7) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(6) => VCC_net_1, MDDR_FABRIC_PWDATA(5)
         => VCC_net_1, MDDR_FABRIC_PWDATA(4) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(3) => VCC_net_1, MDDR_FABRIC_PWDATA(2)
         => VCC_net_1, MDDR_FABRIC_PWDATA(1) => VCC_net_1, 
        MDDR_FABRIC_PWDATA(0) => VCC_net_1, MDDR_FABRIC_PWRITE
         => VCC_net_1, PRESET_N => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => CAN_RX_PAD_Y, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GND_net_1, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => GND_net_1, DM_IN(0) => 
        GND_net_1, DRAM_DQ_IN(17) => GND_net_1, DRAM_DQ_IN(16)
         => GND_net_1, DRAM_DQ_IN(15) => GND_net_1, 
        DRAM_DQ_IN(14) => GND_net_1, DRAM_DQ_IN(13) => GND_net_1, 
        DRAM_DQ_IN(12) => GND_net_1, DRAM_DQ_IN(11) => GND_net_1, 
        DRAM_DQ_IN(10) => GND_net_1, DRAM_DQ_IN(9) => GND_net_1, 
        DRAM_DQ_IN(8) => GND_net_1, DRAM_DQ_IN(7) => GND_net_1, 
        DRAM_DQ_IN(6) => GND_net_1, DRAM_DQ_IN(5) => GND_net_1, 
        DRAM_DQ_IN(4) => GND_net_1, DRAM_DQ_IN(3) => GND_net_1, 
        DRAM_DQ_IN(2) => GND_net_1, DRAM_DQ_IN(1) => GND_net_1, 
        DRAM_DQ_IN(0) => GND_net_1, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => GND_net_1, DRAM_DQS_IN(0) => GND_net_1, 
        DRAM_FIFO_WE_IN(1) => GND_net_1, DRAM_FIFO_WE_IN(0) => 
        GND_net_1, I2C0_SCL_USBC_DATA1_MGPIO31B_IN => 
        I2C_0_SCL_PAD_Y, I2C0_SDA_USBC_DATA0_MGPIO30B_IN => 
        I2C_0_SDA_PAD_Y, I2C1_SCL_USBA_DATA4_MGPIO1A_IN => 
        GPIO_GPIO_1_BI_PAD_Y, I2C1_SDA_USBA_DATA3_MGPIO0A_IN => 
        GND_net_1, MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => 
        GPIO_GPIO_19_BI_PAD_Y, MMUART0_DCD_MGPIO22B_IN => 
        GPIO_GPIO_22_BI_PAD_Y, MMUART0_DSR_MGPIO20B_IN => 
        GPIO_GPIO_20_BI_PAD_Y, MMUART0_DTR_USBC_DATA6_MGPIO18B_IN
         => GND_net_1, MMUART0_RI_MGPIO21B_IN => 
        GPIO_GPIO_21_BI_PAD_Y, MMUART0_RTS_USBC_DATA5_MGPIO17B_IN
         => GND_net_1, MMUART0_RXD_USBC_STP_MGPIO28B_IN => 
        MMUART_0_RXD_PAD_Y, MMUART0_SCK_USBC_NXT_MGPIO29B_IN => 
        GPIO_GPIO_29_BI_PAD_Y, MMUART0_TXD_USBC_DIR_MGPIO27B_IN
         => GND_net_1, MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => 
        GPIO_GPIO_26_BI_PAD_Y, MMUART1_SCK_USBC_DATA4_MGPIO25B_IN
         => GPIO_GPIO_25_BI_PAD_Y, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GPIO_GPIO_8_BI_PAD_Y, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GPIO_GPIO_9_BI_PAD_Y, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GPIO_GPIO_10_BI_PAD_Y, 
        SPI1_SCK_IN => GND_net_1, SPI1_SDI_MGPIO11A_IN => 
        GPIO_GPIO_11_BI_PAD_Y, SPI1_SDO_MGPIO12A_IN => 
        GPIO_GPIO_12_BI_PAD_Y, SPI1_SS0_MGPIO13A_IN => 
        GPIO_GPIO_13_BI_PAD_Y, SPI1_SS1_MGPIO14A_IN => 
        GPIO_GPIO_14_BI_PAD_Y, SPI1_SS2_MGPIO15A_IN => 
        GPIO_GPIO_15_BI_PAD_Y, SPI1_SS3_MGPIO16A_IN => 
        GPIO_GPIO_16_BI_PAD_Y, SPI1_SS4_MGPIO17A_IN => 
        GPIO_GPIO_17_BI_PAD_Y, SPI1_SS5_MGPIO18A_IN => 
        GPIO_GPIO_18_BI_PAD_Y, SPI1_SS6_MGPIO23A_IN => 
        GPIO_GPIO_23_BI_PAD_Y, SPI1_SS7_MGPIO24A_IN => 
        GPIO_GPIO_24_BI_PAD_Y, USBC_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, 
        DRAM_ADDR(15) => nc132, DRAM_ADDR(14) => nc21, 
        DRAM_ADDR(13) => nc237, DRAM_ADDR(12) => nc93, 
        DRAM_ADDR(11) => nc262, DRAM_ADDR(10) => nc69, 
        DRAM_ADDR(9) => nc206, DRAM_ADDR(8) => nc174, 
        DRAM_ADDR(7) => nc38, DRAM_ADDR(6) => nc113, DRAM_ADDR(5)
         => nc218, DRAM_ADDR(4) => nc106, DRAM_ADDR(3) => nc261, 
        DRAM_ADDR(2) => nc25, DRAM_ADDR(1) => nc1, DRAM_ADDR(0)
         => nc299, DRAM_BA(2) => nc37, DRAM_BA(1) => nc202, 
        DRAM_BA(0) => nc144, DRAM_CASN => OPEN, DRAM_CKE => OPEN, 
        DRAM_CLK => OPEN, DRAM_CSN => OPEN, DRAM_DM_RDQS_OUT(2)
         => nc153, DRAM_DM_RDQS_OUT(1) => nc46, 
        DRAM_DM_RDQS_OUT(0) => nc258, DRAM_DQ_OUT(17) => nc71, 
        DRAM_DQ_OUT(16) => nc124, DRAM_DQ_OUT(15) => nc81, 
        DRAM_DQ_OUT(14) => nc201, DRAM_DQ_OUT(13) => nc168, 
        DRAM_DQ_OUT(12) => nc34, DRAM_DQ_OUT(11) => nc28, 
        DRAM_DQ_OUT(10) => nc115, DRAM_DQ_OUT(9) => nc264, 
        DRAM_DQ_OUT(8) => nc192, DRAM_DQ_OUT(7) => nc134, 
        DRAM_DQ_OUT(6) => nc32, DRAM_DQ_OUT(5) => nc40, 
        DRAM_DQ_OUT(4) => nc297, DRAM_DQ_OUT(3) => nc99, 
        DRAM_DQ_OUT(2) => nc75, DRAM_DQ_OUT(1) => nc183, 
        DRAM_DQ_OUT(0) => nc288, DRAM_DQS_OUT(2) => nc85, 
        DRAM_DQS_OUT(1) => nc27, DRAM_DQS_OUT(0) => nc108, 
        DRAM_FIFO_WE_OUT(1) => nc16, DRAM_FIFO_WE_OUT(0) => nc155, 
        DRAM_ODT => OPEN, DRAM_RASN => OPEN, DRAM_RSTN => OPEN, 
        DRAM_WEN => OPEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT => 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT => 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, 
        MMUART0_DCD_MGPIO22B_OUT => 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OUT, 
        MMUART0_DSR_MGPIO20B_OUT => 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OUT, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OUT, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, 
        SPI1_SCK_OUT => OPEN, SPI1_SDI_MGPIO11A_OUT => 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OUT, 
        SPI1_SDO_MGPIO12A_OUT => 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT, 
        SPI1_SS0_MGPIO13A_OUT => 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT, 
        SPI1_SS1_MGPIO14A_OUT => 
        MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OUT, 
        SPI1_SS2_MGPIO15A_OUT => 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OUT, 
        SPI1_SS3_MGPIO16A_OUT => 
        MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OUT, 
        SPI1_SS4_MGPIO17A_OUT => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        SPI1_SS5_MGPIO18A_OUT => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        SPI1_SS6_MGPIO23A_OUT => 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OUT, 
        SPI1_SS7_MGPIO24A_OUT => 
        MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OUT, USBC_XCLK_OUT => 
        OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => OPEN, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => 
        MSS_ADLIB_INST_CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, DM_OE(2)
         => nc51, DM_OE(1) => nc301, DM_OE(0) => nc33, 
        DRAM_DQ_OE(17) => nc204, DRAM_DQ_OE(16) => nc173, 
        DRAM_DQ_OE(15) => nc278, DRAM_DQ_OE(14) => nc169, 
        DRAM_DQ_OE(13) => nc78, DRAM_DQ_OE(12) => nc263, 
        DRAM_DQ_OE(11) => nc24, DRAM_DQ_OE(10) => nc88, 
        DRAM_DQ_OE(9) => nc111, DRAM_DQ_OE(8) => nc55, 
        DRAM_DQ_OE(7) => nc10, DRAM_DQ_OE(6) => nc22, 
        DRAM_DQ_OE(5) => nc210, DRAM_DQ_OE(4) => nc185, 
        DRAM_DQ_OE(3) => nc143, DRAM_DQ_OE(2) => nc248, 
        DRAM_DQ_OE(1) => nc77, DRAM_DQ_OE(0) => nc6, 
        DRAM_DQS_OE(2) => nc109, DRAM_DQS_OE(1) => nc87, 
        DRAM_DQS_OE(0) => nc123, I2C0_SCL_USBC_DATA1_MGPIO31B_OE
         => MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => OPEN, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, 
        MMUART0_DCD_MGPIO22B_OE => 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OE, 
        MMUART0_DSR_MGPIO20B_OE => 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OE, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => 
        MSS_ADLIB_INST_MMUART0_RI_MGPIO21B_OE, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OE, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => 
        MSS_ADLIB_INST_MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => OPEN, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => 
        MSS_ADLIB_INST_SPI0_SS2_USBA_DATA6_MGPIO9A_OE, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OE, 
        SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        MSS_ADLIB_INST_SPI1_SDI_MGPIO11A_OE, SPI1_SDO_MGPIO12A_OE
         => MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE, 
        SPI1_SS0_MGPIO13A_OE => 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE, SPI1_SS1_MGPIO14A_OE
         => MSS_ADLIB_INST_SPI1_SS1_MGPIO14A_OE, 
        SPI1_SS2_MGPIO15A_OE => 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OE, SPI1_SS3_MGPIO16A_OE
         => MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OE, 
        SPI1_SS4_MGPIO17A_OE => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, SPI1_SS5_MGPIO18A_OE
         => MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE => 
        MSS_ADLIB_INST_SPI1_SS6_MGPIO23A_OE, SPI1_SS7_MGPIO24A_OE
         => MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OE, USBC_XCLK_OE => 
        OPEN);
    
    MSS_ADLIB_INST_RNO_5 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(6), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[6]\);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MSS_ADLIB_INST_RNO_25 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(26), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[26]\);
    
    MSS_ADLIB_INST_RNO_24 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(25), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[25]\);
    
    GPIO_GPIO_22_BI_PAD : BIBUF
      port map(PAD => GPIO_22_BI, D => 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_DCD_MGPIO22B_OE, Y => 
        GPIO_GPIO_22_BI_PAD_Y);
    
    GPIO_GPIO_18_BI_PAD : BIBUF
      port map(PAD => GPIO_18_BI, D => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, Y => 
        GPIO_GPIO_18_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_1 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(2), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[2]\);
    
    GPIO_GPIO_16_BI_PAD : BIBUF
      port map(PAD => GPIO_16_BI, D => 
        MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS3_MGPIO16A_OE, Y => 
        GPIO_GPIO_16_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_30 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(31), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[31]\);
    
    I2C_0_SDA_PAD : BIBUF
      port map(PAD => I2C_0_SDA, D => 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, E => 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE, Y => 
        I2C_0_SDA_PAD_Y);
    
    GPIO_GPIO_19_BI_PAD : BIBUF
      port map(PAD => GPIO_19_BI, D => 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, Y => 
        GPIO_GPIO_19_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_26 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(27), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[27]\);
    
    GPIO_GPIO_10_BI_PAD : BIBUF
      port map(PAD => GPIO_10_BI, D => 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS3_USBA_DATA7_MGPIO10A_OE, Y => 
        GPIO_GPIO_10_BI_PAD_Y);
    
    CAN_TX_EN_N_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, E => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, PAD => 
        CAN_TX_EN_N);
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    MSS_ADLIB_INST_RNO_8 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(9), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[9]\);
    
    MSS_ADLIB_INST_RNO_6 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(7), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[7]\);
    
    MSS_ADLIB_INST_RNO_28 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(29), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[29]\);
    
    CAN_RX_PAD : INBUF
      port map(PAD => CAN_RX, Y => CAN_RX_PAD_Y);
    
    GPIO_GPIO_24_BI_PAD : BIBUF
      port map(PAD => GPIO_24_BI, D => 
        MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS7_MGPIO24A_OE, Y => 
        GPIO_GPIO_24_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_9 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(10), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[10]\);
    
    MSS_ADLIB_INST_RNO_15 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(16), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[16]\);
    
    MSS_ADLIB_INST_RNO_0 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(1), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[1]\);
    
    GPIO_GPIO_8_BI_PAD : BIBUF
      port map(PAD => GPIO_8_BI, D => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, Y => 
        GPIO_GPIO_8_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_14 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(15), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[15]\);
    
    GPIO_GPIO_26_BI_PAD : BIBUF
      port map(PAD => GPIO_26_BI, D => 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, Y => 
        GPIO_GPIO_26_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_16 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(17), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[17]\);
    
    GPIO_GPIO_29_BI_PAD : BIBUF
      port map(PAD => GPIO_29_BI, D => 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_SCK_USBC_NXT_MGPIO29B_OE, Y => 
        GPIO_GPIO_29_BI_PAD_Y);
    
    GPIO_GPIO_20_BI_PAD : BIBUF
      port map(PAD => GPIO_20_BI, D => 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OUT, E => 
        MSS_ADLIB_INST_MMUART0_DSR_MGPIO20B_OE, Y => 
        GPIO_GPIO_20_BI_PAD_Y);
    
    GPIO_GPIO_15_BI_PAD : BIBUF
      port map(PAD => GPIO_15_BI, D => 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS2_MGPIO15A_OE, Y => 
        GPIO_GPIO_15_BI_PAD_Y);
    
    MSS_ADLIB_INST_RNO_18 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(19), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[19]\);
    
    MSS_ADLIB_INST_RNO_3 : CFG2
      generic map(INIT => x"8")

      port map(A => hready_m_xhdl349, B => 
        CoreAHBLite_0_AHBmslave10_HRDATA(4), Y => 
        \CoreAHBLite_0_AHBmslave10_HRDATA_m[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_slave_stage is

    port( AWSIZE_IS16_gated               : in    std_logic_vector(1 downto 0);
          ARADDR_IS16_gated               : in    std_logic_vector(23 downto 1);
          AWADDR_IS16_gated               : in    std_logic_vector(23 downto 1);
          ARSIZE_IS16_gated               : in    std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_ARSIZE    : out   std_logic_vector(1 downto 0);
          WDATA_IS16_gated                : in    std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_WDATA     : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated                : in    std_logic_vector(7 downto 0);
          COREAXI_0_AXImslave16_WSTRB     : out   std_logic_vector(7 downto 0);
          COREAXI_0_AXImslave16_AWADDR    : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_ARADDR    : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_AWSIZE    : out   std_logic_vector(1 downto 0);
          ARBURST_IS16_gated_0            : in    std_logic;
          COREAXI_0_AXImslave16_ARBURST_0 : out   std_logic;
          WREADY_SI16                     : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY   : in    std_logic;
          COREAXI_0_AXImslave16_AWREADY   : in    std_logic;
          WVALID_IS16                     : in    std_logic;
          AWVALID_IS16                    : in    std_logic;
          ARVALID_IS16                    : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID   : out   std_logic;
          AWREADY_SI16                    : out   std_logic;
          COREAXI_0_AXImslave16_AWVALID   : out   std_logic;
          WREADY_SI16_i                   : in    std_logic;
          COREAXI_0_AXImslave16_WVALID    : out   std_logic;
          SDRCLK_c                        : in    std_logic;
          MSS_READY                       : in    std_logic
        );

end axi_slave_stage;

architecture DEF_ARCH of axi_slave_stage is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_2755_i, \AWVALID_S_xhdl20_1_sqmuxa_i\, 
        GND_net_1, N_2743_i, N_2731_i, 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, N_2720_i, N_2709_i, 
        N_2698_i, N_2687_i, N_2676_i, N_2665_i, N_2654_i, 
        N_2643_i, N_2632_i, N_2621_i, N_2530_i, N_2519_i, 
        N_2508_i, N_2497_i, N_2486_i, N_2475_i, N_2464_i, 
        N_2453_i, N_2442_i, N_2431_i, N_2420_i, N_2409_i, 
        N_2398_i, N_2386_i, N_2374_i, N_2362_i, N_2350_i, 
        N_2338_i, N_2326_i, N_2314_i, N_2302_i, N_2290_i, 
        N_2218_i, N_2206_i, N_2194_i, N_2182_i, N_2170_i, 
        N_2158_i, N_2146_i, N_2134_i, N_2122_i, N_2110_i, 
        N_2098_i, N_2086_i, N_2074_i, N_3162_i, N_2062_i, 
        N_2051_i, N_2016_i, \WLAST_S_xhdl24_1_sqmuxa_i_0\, 
        \COREAXI_0_AXImslave16_AWVALID\, \AWREADY_SI16\, 
        \COREAXI_0_AXImslave16_ARVALID\, ARREADY_SI16_i, 
        \ARVALID_IS_r\, \AWVALID_IS_r\, \WVALID_IS_r\, 
        \AWVALID_IS_r1\, \WVALID_IS_r1\ : std_logic;

begin 

    COREAXI_0_AXImslave16_ARVALID <= 
        \COREAXI_0_AXImslave16_ARVALID\;
    AWREADY_SI16 <= \AWREADY_SI16\;
    COREAXI_0_AXImslave16_AWVALID <= 
        \COREAXI_0_AXImslave16_AWVALID\;

    \ARADDR_S_xhdl28_RNO[5]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(5), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2486_i);
    
    ARVALID_S_xhdl35_1_sqmuxa_i : CFG4
      generic map(INIT => x"AE0C")

      port map(A => \COREAXI_0_AXImslave16_ARVALID\, B => 
        ARVALID_IS16, C => \ARVALID_IS_r\, D => 
        COREAXI_0_AXImslave16_ARREADY, Y => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\);
    
    \WDATA_S_xhdl22[56]\ : SLE
      port map(D => WDATA_IS16_gated(56), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(56));
    
    \AWADDR_S_xhdl13_RNO[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(6), Y
         => N_2158_i);
    
    \ARADDR_S_xhdl28[19]\ : SLE
      port map(D => N_2665_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(19));
    
    \ARADDR_S_xhdl28[18]\ : SLE
      port map(D => N_2676_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(18));
    
    \ARADDR_S_xhdl28[8]\ : SLE
      port map(D => N_2453_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(8));
    
    \AWADDR_S_xhdl13_RNO[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(8), Y
         => N_2134_i);
    
    \WSTRB_S_xhdl23[4]\ : SLE
      port map(D => WSTRB_IS16_gated(4), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(4));
    
    \ARSIZE_S_xhdl30_RNO[1]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARSIZE_IS16_gated(1), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2051_i);
    
    \WSTRB_S_xhdl23[7]\ : SLE
      port map(D => WSTRB_IS16_gated(7), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(7));
    
    \AWADDR_S_xhdl13_RNO[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(15), Y
         => N_2386_i);
    
    AWVALID_S_xhdl20_1_sqmuxa_i : CFG4
      generic map(INIT => x"10FF")

      port map(A => \AWVALID_IS_r1\, B => \AWVALID_IS_r\, C => 
        AWVALID_IS16, D => \AWREADY_SI16\, Y => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\);
    
    \WDATA_S_xhdl22[40]\ : SLE
      port map(D => WDATA_IS16_gated(40), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(40));
    
    \WDATA_S_xhdl22[30]\ : SLE
      port map(D => WDATA_IS16_gated(30), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(30));
    
    \ARADDR_S_xhdl28_RNO[21]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(21), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2643_i);
    
    \ARADDR_S_xhdl28_RNO[13]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(13), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2731_i);
    
    \ARADDR_S_xhdl28_RNO[10]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(10), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2431_i);
    
    \WDATA_S_xhdl22[50]\ : SLE
      port map(D => WDATA_IS16_gated(50), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(50));
    
    \WDATA_S_xhdl22[49]\ : SLE
      port map(D => WDATA_IS16_gated(49), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(49));
    
    \WDATA_S_xhdl22[39]\ : SLE
      port map(D => WDATA_IS16_gated(39), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(39));
    
    \WDATA_S_xhdl22[47]\ : SLE
      port map(D => WDATA_IS16_gated(47), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(47));
    
    \WDATA_S_xhdl22[37]\ : SLE
      port map(D => WDATA_IS16_gated(37), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(37));
    
    \AWSIZE_S_xhdl15[1]\ : SLE
      port map(D => N_2743_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWSIZE(1));
    
    \WDATA_S_xhdl22[18]\ : SLE
      port map(D => WDATA_IS16_gated(18), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(18));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \AWADDR_S_xhdl13[21]\ : SLE
      port map(D => N_2314_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(21));
    
    \WDATA_S_xhdl22[59]\ : SLE
      port map(D => WDATA_IS16_gated(59), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(59));
    
    \WDATA_S_xhdl22[57]\ : SLE
      port map(D => WDATA_IS16_gated(57), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(57));
    
    \AWADDR_S_xhdl13[8]\ : SLE
      port map(D => N_2134_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(8));
    
    \AWADDR_S_xhdl13[17]\ : SLE
      port map(D => N_2362_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(17));
    
    \ARADDR_S_xhdl28_RNO[8]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(8), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2453_i);
    
    \ARADDR_S_xhdl28_RNO[6]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(6), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2475_i);
    
    \AWADDR_S_xhdl13[10]\ : SLE
      port map(D => N_2110_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(10));
    
    ARVALID_S_xhdl35 : SLE
      port map(D => ARREADY_SI16_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \COREAXI_0_AXImslave16_ARVALID\);
    
    \AWADDR_S_xhdl13[1]\ : SLE
      port map(D => N_2218_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(1));
    
    \WDATA_S_xhdl22[16]\ : SLE
      port map(D => WDATA_IS16_gated(16), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(16));
    
    \WDATA_S_xhdl22[41]\ : SLE
      port map(D => WDATA_IS16_gated(41), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(41));
    
    \WDATA_S_xhdl22[31]\ : SLE
      port map(D => WDATA_IS16_gated(31), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(31));
    
    \AWADDR_S_xhdl13_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(1), Y
         => N_2218_i);
    
    \WDATA_S_xhdl22[28]\ : SLE
      port map(D => WDATA_IS16_gated(28), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(28));
    
    \WDATA_S_xhdl22[42]\ : SLE
      port map(D => WDATA_IS16_gated(42), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(42));
    
    \WDATA_S_xhdl22[32]\ : SLE
      port map(D => WDATA_IS16_gated(32), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(32));
    
    \ARADDR_S_xhdl28_RNO[17]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(17), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2687_i);
    
    \WSTRB_S_xhdl23[0]\ : SLE
      port map(D => WSTRB_IS16_gated(0), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(0));
    
    \WDATA_S_xhdl22[51]\ : SLE
      port map(D => WDATA_IS16_gated(51), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(51));
    
    \WDATA_S_xhdl22[44]\ : SLE
      port map(D => WDATA_IS16_gated(44), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(44));
    
    \WDATA_S_xhdl22[34]\ : SLE
      port map(D => WDATA_IS16_gated(34), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(34));
    
    \WDATA_S_xhdl22[52]\ : SLE
      port map(D => WDATA_IS16_gated(52), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(52));
    
    \AWADDR_S_xhdl13_RNO[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(16), Y
         => N_2374_i);
    
    ARVALID_IS_r : SLE
      port map(D => ARVALID_IS16, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARVALID_IS_r\);
    
    \WSTRB_S_xhdl23[5]\ : SLE
      port map(D => WSTRB_IS16_gated(5), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(5));
    
    \ARADDR_S_xhdl28_RNO[12]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(12), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2409_i);
    
    \WDATA_S_xhdl22[54]\ : SLE
      port map(D => WDATA_IS16_gated(54), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(54));
    
    \WDATA_S_xhdl22[26]\ : SLE
      port map(D => WDATA_IS16_gated(26), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(26));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \AWADDR_S_xhdl13[12]\ : SLE
      port map(D => N_2086_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(12));
    
    \WDATA_S_xhdl22[7]\ : SLE
      port map(D => WDATA_IS16_gated(7), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(7));
    
    \AWADDR_S_xhdl13_RNO[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(4), Y
         => N_2182_i);
    
    \AWSIZE_S_xhdl15_RNO[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWSIZE_IS16_gated(0), Y
         => N_2755_i);
    
    \AWADDR_S_xhdl13_RNO[17]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(17), Y
         => N_2362_i);
    
    \ARADDR_S_xhdl28_RNO[16]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(16), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2698_i);
    
    \AWADDR_S_xhdl13_RNO[23]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(23), Y
         => N_2290_i);
    
    \WDATA_S_xhdl22[10]\ : SLE
      port map(D => WDATA_IS16_gated(10), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(10));
    
    \ARADDR_S_xhdl28_RNO[2]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(2), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2519_i);
    
    \WDATA_S_xhdl22[0]\ : SLE
      port map(D => WDATA_IS16_gated(0), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(0));
    
    \AWADDR_S_xhdl13[23]\ : SLE
      port map(D => N_2290_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(23));
    
    AWVALID_IS_r : SLE
      port map(D => AWVALID_IS16, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWVALID_IS_r\);
    
    \AWADDR_S_xhdl13_RNO[22]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(22), Y
         => N_2302_i);
    
    WVALID_IS_r : SLE
      port map(D => WVALID_IS16, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \WVALID_IS_r\);
    
    WLAST_S_xhdl24_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"FF10")

      port map(A => \WVALID_IS_r1\, B => \WVALID_IS_r\, C => 
        WVALID_IS16, D => WREADY_SI16, Y => 
        \WLAST_S_xhdl24_1_sqmuxa_i_0\);
    
    \ARADDR_S_xhdl28[15]\ : SLE
      port map(D => N_2709_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(15));
    
    \WDATA_S_xhdl22[19]\ : SLE
      port map(D => WDATA_IS16_gated(19), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(19));
    
    \AWADDR_S_xhdl13_RNO[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(20), Y
         => N_2326_i);
    
    \WDATA_S_xhdl22[17]\ : SLE
      port map(D => WDATA_IS16_gated(17), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(17));
    
    \WDATA_S_xhdl22[60]\ : SLE
      port map(D => WDATA_IS16_gated(60), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(60));
    
    \AWADDR_S_xhdl13_RNO[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(7), Y
         => N_2146_i);
    
    AWVALID_S_xhdl20 : SLE
      port map(D => \AWREADY_SI16\, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \COREAXI_0_AXImslave16_AWVALID\);
    
    \AWSIZE_S_xhdl15[0]\ : SLE
      port map(D => N_2755_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWSIZE(0));
    
    \AWADDR_S_xhdl13_RNO[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(2), Y
         => N_2206_i);
    
    \AWADDR_S_xhdl13_RNO[19]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(19), Y
         => N_2338_i);
    
    \WDATA_S_xhdl22[20]\ : SLE
      port map(D => WDATA_IS16_gated(20), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(20));
    
    \AWADDR_S_xhdl13[15]\ : SLE
      port map(D => N_2386_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(15));
    
    \WDATA_S_xhdl22[43]\ : SLE
      port map(D => WDATA_IS16_gated(43), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(43));
    
    \WDATA_S_xhdl22[33]\ : SLE
      port map(D => WDATA_IS16_gated(33), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(33));
    
    \AWADDR_S_xhdl13[4]\ : SLE
      port map(D => N_2182_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(4));
    
    \WDATA_S_xhdl22[29]\ : SLE
      port map(D => WDATA_IS16_gated(29), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(29));
    
    AWVALID_IS_r1 : SLE
      port map(D => \AWVALID_IS_r\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWVALID_IS_r1\);
    
    \AWADDR_S_xhdl13_RNO[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(3), Y
         => N_2194_i);
    
    \WDATA_S_xhdl22[27]\ : SLE
      port map(D => WDATA_IS16_gated(27), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(27));
    
    \WDATA_S_xhdl22[11]\ : SLE
      port map(D => WDATA_IS16_gated(11), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(11));
    
    \AWADDR_S_xhdl13[18]\ : SLE
      port map(D => N_2350_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(18));
    
    \ARADDR_S_xhdl28[21]\ : SLE
      port map(D => N_2643_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(21));
    
    \WDATA_S_xhdl22[4]\ : SLE
      port map(D => WDATA_IS16_gated(4), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(4));
    
    \WDATA_S_xhdl22[12]\ : SLE
      port map(D => WDATA_IS16_gated(12), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(12));
    
    AWREADY_SI : CFG2
      generic map(INIT => x"7")

      port map(A => \COREAXI_0_AXImslave16_AWVALID\, B => 
        COREAXI_0_AXImslave16_AWREADY, Y => \AWREADY_SI16\);
    
    \ARADDR_S_xhdl28[11]\ : SLE
      port map(D => N_2420_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(11));
    
    \WDATA_S_xhdl22[53]\ : SLE
      port map(D => WDATA_IS16_gated(53), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(53));
    
    \AWSIZE_S_xhdl15_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWSIZE_IS16_gated(1), Y
         => N_2743_i);
    
    \AWADDR_S_xhdl13_RNO[14]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(14), Y
         => N_2398_i);
    
    \WSTRB_S_xhdl23[6]\ : SLE
      port map(D => WSTRB_IS16_gated(6), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(6));
    
    \ARADDR_S_xhdl28[22]\ : SLE
      port map(D => N_2632_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(22));
    
    \WDATA_S_xhdl22[14]\ : SLE
      port map(D => WDATA_IS16_gated(14), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(14));
    
    \AWADDR_S_xhdl13[7]\ : SLE
      port map(D => N_2146_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(7));
    
    \ARADDR_S_xhdl28[12]\ : SLE
      port map(D => N_2409_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(12));
    
    \WDATA_S_xhdl22[61]\ : SLE
      port map(D => WDATA_IS16_gated(61), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(61));
    
    \ARADDR_S_xhdl28_RNO[11]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(11), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2420_i);
    
    \WDATA_S_xhdl22[45]\ : SLE
      port map(D => WDATA_IS16_gated(45), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(45));
    
    \WDATA_S_xhdl22[35]\ : SLE
      port map(D => WDATA_IS16_gated(35), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(35));
    
    \WDATA_S_xhdl22[1]\ : SLE
      port map(D => WDATA_IS16_gated(1), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(1));
    
    \AWADDR_S_xhdl13_RNO[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(9), Y
         => N_2122_i);
    
    \WDATA_S_xhdl22[62]\ : SLE
      port map(D => WDATA_IS16_gated(62), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(62));
    
    \AWADDR_S_xhdl13_RNO[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(13), Y
         => N_2074_i);
    
    \ARADDR_S_xhdl28_RNO[4]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(4), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2497_i);
    
    \WDATA_S_xhdl22[9]\ : SLE
      port map(D => WDATA_IS16_gated(9), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(9));
    
    \WDATA_S_xhdl22[21]\ : SLE
      port map(D => WDATA_IS16_gated(21), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(21));
    
    \WDATA_S_xhdl22[55]\ : SLE
      port map(D => WDATA_IS16_gated(55), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(55));
    
    \AWADDR_S_xhdl13[11]\ : SLE
      port map(D => N_2098_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(11));
    
    \WDATA_S_xhdl22[22]\ : SLE
      port map(D => WDATA_IS16_gated(22), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(22));
    
    \AWADDR_S_xhdl13[19]\ : SLE
      port map(D => N_2338_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(19));
    
    \AWADDR_S_xhdl13_RNO[12]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(12), Y
         => N_2086_i);
    
    \ARADDR_S_xhdl28_RNO[19]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(19), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2665_i);
    
    \AWADDR_S_xhdl13_RNO[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(21), Y
         => N_2314_i);
    
    \ARBURST_S_xhdl31_RNO[0]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARBURST_IS16_gated_0, B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2016_i);
    
    \AWADDR_S_xhdl13_RNO[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(10), Y
         => N_2110_i);
    
    \ARADDR_S_xhdl28_RNO[23]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(23), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2621_i);
    
    \ARADDR_S_xhdl28_RNO[20]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(20), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2654_i);
    
    WVALID_IS_r1 : SLE
      port map(D => \WVALID_IS_r\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WVALID_IS_r1\);
    
    \WDATA_S_xhdl22[24]\ : SLE
      port map(D => WDATA_IS16_gated(24), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(24));
    
    \WDATA_S_xhdl22[6]\ : SLE
      port map(D => WDATA_IS16_gated(6), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(6));
    
    \ARSIZE_S_xhdl30[0]\ : SLE
      port map(D => N_2062_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARSIZE(0));
    
    \WSTRB_S_xhdl23[1]\ : SLE
      port map(D => WSTRB_IS16_gated(1), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(1));
    
    \ARBURST_S_xhdl31[0]\ : SLE
      port map(D => N_2016_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARBURST_0);
    
    \ARADDR_S_xhdl28[14]\ : SLE
      port map(D => N_2720_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(14));
    
    \WDATA_S_xhdl22[5]\ : SLE
      port map(D => WDATA_IS16_gated(5), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(5));
    
    \ARADDR_S_xhdl28[2]\ : SLE
      port map(D => N_2519_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(2));
    
    \WDATA_S_xhdl22[3]\ : SLE
      port map(D => WDATA_IS16_gated(3), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(3));
    
    \ARADDR_S_xhdl28[20]\ : SLE
      port map(D => N_2654_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(20));
    
    WVALID_IS_r1_RNI619R : CFG4
      generic map(INIT => x"0010")

      port map(A => \WVALID_IS_r1\, B => \WVALID_IS_r\, C => 
        WVALID_IS16, D => WREADY_SI16, Y => N_3162_i);
    
    \ARADDR_S_xhdl28[10]\ : SLE
      port map(D => N_2431_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(10));
    
    \WSTRB_S_xhdl23[3]\ : SLE
      port map(D => WSTRB_IS16_gated(3), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(3));
    
    \ARADDR_S_xhdl28_RNO[9]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(9), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2442_i);
    
    \AWADDR_S_xhdl13[14]\ : SLE
      port map(D => N_2398_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(14));
    
    \WDATA_S_xhdl22[2]\ : SLE
      port map(D => WDATA_IS16_gated(2), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(2));
    
    \ARADDR_S_xhdl28_RNO[15]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(15), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2709_i);
    
    \ARSIZE_S_xhdl30[1]\ : SLE
      port map(D => N_2051_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARSIZE(1));
    
    \WDATA_S_xhdl22[8]\ : SLE
      port map(D => WDATA_IS16_gated(8), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(8));
    
    \AWADDR_S_xhdl13[20]\ : SLE
      port map(D => N_2326_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(20));
    
    \ARADDR_S_xhdl28[6]\ : SLE
      port map(D => N_2475_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(6));
    
    ARVALID_S_xhdl35_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => \COREAXI_0_AXImslave16_ARVALID\, B => 
        COREAXI_0_AXImslave16_ARREADY, Y => ARREADY_SI16_i);
    
    \ARADDR_S_xhdl28[3]\ : SLE
      port map(D => N_2508_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(3));
    
    \AWADDR_S_xhdl13[2]\ : SLE
      port map(D => N_2206_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(2));
    
    \ARADDR_S_xhdl28_RNO[18]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(18), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2676_i);
    
    \WDATA_S_xhdl22[13]\ : SLE
      port map(D => WDATA_IS16_gated(13), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(13));
    
    \ARADDR_S_xhdl28_RNO[14]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(14), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2720_i);
    
    \AWADDR_S_xhdl13[16]\ : SLE
      port map(D => N_2374_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(16));
    
    \ARADDR_S_xhdl28[7]\ : SLE
      port map(D => N_2464_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(7));
    
    \ARADDR_S_xhdl28[16]\ : SLE
      port map(D => N_2698_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(16));
    
    \ARADDR_S_xhdl28[1]\ : SLE
      port map(D => N_2530_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(1));
    
    \ARADDR_S_xhdl28_RNO[7]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(7), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2464_i);
    
    \ARADDR_S_xhdl28[23]\ : SLE
      port map(D => N_2621_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(23));
    
    \WDATA_S_xhdl22[63]\ : SLE
      port map(D => WDATA_IS16_gated(63), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(63));
    
    \AWADDR_S_xhdl13[6]\ : SLE
      port map(D => N_2158_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(6));
    
    \AWADDR_S_xhdl13[13]\ : SLE
      port map(D => N_2074_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(13));
    
    \ARADDR_S_xhdl28_RNO[22]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(22), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2632_i);
    
    \ARADDR_S_xhdl28[13]\ : SLE
      port map(D => N_2731_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(13));
    
    \WSTRB_S_xhdl23[2]\ : SLE
      port map(D => WSTRB_IS16_gated(2), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WSTRB(2));
    
    \WDATA_S_xhdl22[15]\ : SLE
      port map(D => WDATA_IS16_gated(15), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(15));
    
    \WDATA_S_xhdl22[48]\ : SLE
      port map(D => WDATA_IS16_gated(48), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(48));
    
    \WDATA_S_xhdl22[38]\ : SLE
      port map(D => WDATA_IS16_gated(38), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(38));
    
    \AWADDR_S_xhdl13_RNO[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(11), Y
         => N_2098_i);
    
    \ARSIZE_S_xhdl30_RNO[0]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARSIZE_IS16_gated(0), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2062_i);
    
    WVALID_S_xhdl25 : SLE
      port map(D => WREADY_SI16_i, CLK => SDRCLK_c, EN => 
        \WLAST_S_xhdl24_1_sqmuxa_i_0\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_WVALID);
    
    \WDATA_S_xhdl22[23]\ : SLE
      port map(D => WDATA_IS16_gated(23), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(23));
    
    \AWADDR_S_xhdl13[22]\ : SLE
      port map(D => N_2302_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(22));
    
    \WDATA_S_xhdl22[58]\ : SLE
      port map(D => WDATA_IS16_gated(58), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(58));
    
    \ARADDR_S_xhdl28[4]\ : SLE
      port map(D => N_2497_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(4));
    
    \ARADDR_S_xhdl28[17]\ : SLE
      port map(D => N_2687_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(17));
    
    \AWADDR_S_xhdl13_RNO[18]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(18), Y
         => N_2350_i);
    
    \AWADDR_S_xhdl13[3]\ : SLE
      port map(D => N_2194_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(3));
    
    \AWADDR_S_xhdl13_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \AWREADY_SI16\, B => AWADDR_IS16_gated(5), Y
         => N_2170_i);
    
    \WDATA_S_xhdl22[46]\ : SLE
      port map(D => WDATA_IS16_gated(46), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(46));
    
    \WDATA_S_xhdl22[36]\ : SLE
      port map(D => WDATA_IS16_gated(36), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(36));
    
    \WDATA_S_xhdl22[25]\ : SLE
      port map(D => WDATA_IS16_gated(25), CLK => SDRCLK_c, EN => 
        N_3162_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAXI_0_AXImslave16_WDATA(25));
    
    \ARADDR_S_xhdl28_RNO[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(3), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2508_i);
    
    \ARADDR_S_xhdl28[9]\ : SLE
      port map(D => N_2442_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(9));
    
    \AWADDR_S_xhdl13[9]\ : SLE
      port map(D => N_2122_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(9));
    
    \ARADDR_S_xhdl28_RNO[1]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => ARADDR_IS16_gated(1), B => 
        COREAXI_0_AXImslave16_ARREADY, C => 
        \COREAXI_0_AXImslave16_ARVALID\, Y => N_2530_i);
    
    \AWADDR_S_xhdl13[5]\ : SLE
      port map(D => N_2170_i, CLK => SDRCLK_c, EN => 
        \AWVALID_S_xhdl20_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_AWADDR(5));
    
    \ARADDR_S_xhdl28[5]\ : SLE
      port map(D => N_2486_i, CLK => SDRCLK_c, EN => 
        \ARVALID_S_xhdl35_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => COREAXI_0_AXImslave16_ARADDR(5));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_master_stage is

    port( RDATA_IM0                            : in    std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : in    std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : in    std_logic_vector(27 downto 1);
          AWADDR_MI0                           : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : out   std_logic_vector(27 downto 1);
          ARSIZE_MI0                           : out   std_logic_vector(1 downto 0);
          AWSIZE_MI0                           : out   std_logic_vector(1 downto 0);
          WDATA_MI0                            : out   std_logic_vector(63 downto 0);
          WSTRB_MI0                            : out   std_logic_vector(7 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : in    std_logic_vector(63 downto 16);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : out   std_logic_vector(63 downto 0);
          axi_current_state_0                  : in    std_logic;
          axi_current_state_3                  : in    std_logic;
          ARBURST_MI0_0                        : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          AWLOCK_MI0_i_0                       : out   std_logic;
          ARLOCK_MI0_i_0                       : out   std_logic;
          ARREADY_IM0                          : in    std_logic;
          awaddr_awvalid_clr_d                 : in    std_logic;
          RVALID_IM0                           : in    std_logic;
          RLAST_IM0                            : in    std_logic;
          AWREADY_IM0                          : in    std_logic;
          WREADY_IM0                           : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : in    std_logic;
          RREADY_MI0                           : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic;
          araddr_arvalid_clr_d                 : in    std_logic;
          BVALID_IM0                           : in    std_logic;
          m0_rd_end                            : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : out   std_logic;
          m0_wr_end                            : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : out   std_logic;
          WVALID_MI0                           : out   std_logic;
          N_48                                 : in    std_logic;
          AWVALID_MI0                          : out   std_logic;
          ARVALID_MI0                          : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          N_75_i                               : in    std_logic;
          N_135_i                              : in    std_logic;
          N_136_i                              : in    std_logic;
          N_137_i                              : in    std_logic;
          N_203_i                              : in    std_logic;
          N_272_i                              : in    std_logic;
          N_273_i                              : in    std_logic;
          N_274_i                              : in    std_logic;
          N_275_i                              : in    std_logic;
          N_276_i                              : in    std_logic;
          N_277_i                              : in    std_logic;
          N_382_i                              : in    std_logic;
          N_381_i                              : in    std_logic;
          N_278_i                              : in    std_logic;
          N_380_i                              : in    std_logic;
          N_133_i                              : in    std_logic;
          N_134_i                              : in    std_logic;
          N_195_i                              : in    std_logic;
          N_197_i                              : in    std_logic;
          N_200_i                              : in    std_logic;
          N_201_i                              : in    std_logic;
          N_202_i                              : in    std_logic;
          N_1452_i                             : in    std_logic;
          N_1451_i                             : in    std_logic;
          N_1450_i                             : in    std_logic;
          N_1449_i                             : in    std_logic;
          N_1448_i                             : in    std_logic;
          N_1447_i                             : in    std_logic;
          N_1446_i                             : in    std_logic;
          N_1445_i                             : in    std_logic;
          wready_m_xhdl2                       : out   std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : out   std_logic
        );

end axi_master_stage;

architecture DEF_ARCH of axi_master_stage is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID_i, 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY_i, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY_i, \ARLOCK_MI0[1]\, 
        \AWLOCK_MI0[1]\, VCC_net_1, \RDATA_M_xhdl8_3[49]\, 
        GND_net_1, \RDATA_M_xhdl8_3[50]\, \RDATA_M_xhdl8_3[51]\, 
        \RDATA_M_xhdl8_3[52]\, \RDATA_M_xhdl8_3[53]\, 
        \RDATA_M_xhdl8_3[54]\, \RDATA_M_xhdl8_3[55]\, 
        \RDATA_M_xhdl8_3[56]\, \RDATA_M_xhdl8_3[57]\, 
        \RDATA_M_xhdl8_3[58]\, \RDATA_M_xhdl8_3[59]\, 
        \RDATA_M_xhdl8_3[60]\, \RDATA_M_xhdl8_3[61]\, 
        \RDATA_M_xhdl8_3[62]\, \RDATA_M_xhdl8_3[63]\, 
        \RDATA_M_xhdl8_3[34]\, \RDATA_M_xhdl8_3[35]\, 
        \RDATA_M_xhdl8_3[36]\, \RDATA_M_xhdl8_3[37]\, 
        \RDATA_M_xhdl8_3[38]\, \RDATA_M_xhdl8_3[39]\, 
        \RDATA_M_xhdl8_3[40]\, \RDATA_M_xhdl8_3[41]\, 
        \RDATA_M_xhdl8_3[42]\, \RDATA_M_xhdl8_3[43]\, 
        \RDATA_M_xhdl8_3[44]\, \RDATA_M_xhdl8_3[45]\, 
        \RDATA_M_xhdl8_3[46]\, \RDATA_M_xhdl8_3[47]\, 
        \RDATA_M_xhdl8_3[48]\, \RDATA_M_xhdl8_3[19]\, 
        \RDATA_M_xhdl8_3[20]\, \RDATA_M_xhdl8_3[21]\, 
        \RDATA_M_xhdl8_3[22]\, \RDATA_M_xhdl8_3[23]\, 
        \RDATA_M_xhdl8_3[24]\, \RDATA_M_xhdl8_3[25]\, 
        \RDATA_M_xhdl8_3[26]\, \RDATA_M_xhdl8_3[27]\, 
        \RDATA_M_xhdl8_3[28]\, \RDATA_M_xhdl8_3[29]\, 
        \RDATA_M_xhdl8_3[30]\, \RDATA_M_xhdl8_3[31]\, 
        \RDATA_M_xhdl8_3[32]\, \RDATA_M_xhdl8_3[33]\, 
        \RDATA_M_xhdl8_3[4]\, \RDATA_M_xhdl8_3[5]\, 
        \RDATA_M_xhdl8_3[6]\, \RDATA_M_xhdl8_3[7]\, 
        \RDATA_M_xhdl8_3[8]\, \RDATA_M_xhdl8_3[9]\, 
        \RDATA_M_xhdl8_3[10]\, \RDATA_M_xhdl8_3[11]\, 
        \RDATA_M_xhdl8_3[12]\, \RDATA_M_xhdl8_3[13]\, 
        \RDATA_M_xhdl8_3[14]\, \RDATA_M_xhdl8_3[15]\, 
        \RDATA_M_xhdl8_3[16]\, \RDATA_M_xhdl8_3[17]\, 
        \RDATA_M_xhdl8_3[18]\, \rd_wdcntr[0]_net_1\, N_16_i, 
        \rd_wdcntr[1]_net_1\, N_22_i, \rd_wdcntr[2]_net_1\, 
        N_20_i, \rd_wdcntr[3]_net_1\, N_18_i, 
        \RDATA_M_xhdl8_3[0]\, \RDATA_M_xhdl8_3[1]\, 
        \RDATA_M_xhdl8_3[2]\, \RDATA_M_xhdl8_3[3]\, 
        \RDATA_M_int[63]_net_1\, \RDATA_M_int_2[63]\, 
        \RDATA_M_int[48]_net_1\, \RDATA_M_int_2[48]\, 
        \RDATA_M_int[49]_net_1\, \RDATA_M_int_2[49]\, 
        \RDATA_M_int[50]_net_1\, \RDATA_M_int_2[50]\, 
        \RDATA_M_int[51]_net_1\, \RDATA_M_int_2[51]\, 
        \RDATA_M_int[52]_net_1\, \RDATA_M_int_2[52]\, 
        \RDATA_M_int[53]_net_1\, \RDATA_M_int_2[53]\, 
        \RDATA_M_int[54]_net_1\, \RDATA_M_int_2[54]\, 
        \RDATA_M_int[55]_net_1\, \RDATA_M_int_2[55]\, 
        \RDATA_M_int[56]_net_1\, \RDATA_M_int_2[56]\, 
        \RDATA_M_int[57]_net_1\, \RDATA_M_int_2[57]\, 
        \RDATA_M_int[58]_net_1\, \RDATA_M_int_2[58]\, 
        \RDATA_M_int[59]_net_1\, \RDATA_M_int_2[59]\, 
        \RDATA_M_int[60]_net_1\, \RDATA_M_int_2[60]\, 
        \RDATA_M_int[61]_net_1\, \RDATA_M_int_2[61]\, 
        \RDATA_M_int[62]_net_1\, \RDATA_M_int_2[62]\, 
        \RDATA_M_int[33]_net_1\, \RDATA_M_int_2[33]\, 
        \RDATA_M_int[34]_net_1\, \RDATA_M_int_2[34]\, 
        \RDATA_M_int[35]_net_1\, \RDATA_M_int_2[35]\, 
        \RDATA_M_int[36]_net_1\, \RDATA_M_int_2[36]\, 
        \RDATA_M_int[37]_net_1\, \RDATA_M_int_2[37]\, 
        \RDATA_M_int[38]_net_1\, \RDATA_M_int_2[38]\, 
        \RDATA_M_int[39]_net_1\, \RDATA_M_int_2[39]\, 
        \RDATA_M_int[40]_net_1\, \RDATA_M_int_2[40]\, 
        \RDATA_M_int[41]_net_1\, \RDATA_M_int_2[41]\, 
        \RDATA_M_int[42]_net_1\, \RDATA_M_int_2[42]\, 
        \RDATA_M_int[43]_net_1\, \RDATA_M_int_2[43]\, 
        \RDATA_M_int[44]_net_1\, \RDATA_M_int_2[44]\, 
        \RDATA_M_int[45]_net_1\, \RDATA_M_int_2[45]\, 
        \RDATA_M_int[46]_net_1\, \RDATA_M_int_2[46]\, 
        \RDATA_M_int[47]_net_1\, \RDATA_M_int_2[47]\, 
        \RDATA_M_int[18]_net_1\, \RDATA_M_int_2[18]\, 
        \RDATA_M_int[19]_net_1\, \RDATA_M_int_2[19]\, 
        \RDATA_M_int[20]_net_1\, \RDATA_M_int_2[20]\, 
        \RDATA_M_int[21]_net_1\, \RDATA_M_int_2[21]\, 
        \RDATA_M_int[22]_net_1\, \RDATA_M_int_2[22]\, 
        \RDATA_M_int[23]_net_1\, \RDATA_M_int_2[23]\, 
        \RDATA_M_int[24]_net_1\, \RDATA_M_int_2[24]\, 
        \RDATA_M_int[25]_net_1\, \RDATA_M_int_2[25]\, 
        \RDATA_M_int[26]_net_1\, \RDATA_M_int_2[26]\, 
        \RDATA_M_int[27]_net_1\, \RDATA_M_int_2[27]\, 
        \RDATA_M_int[28]_net_1\, \RDATA_M_int_2[28]\, 
        \RDATA_M_int[29]_net_1\, \RDATA_M_int_2[29]\, 
        \RDATA_M_int[30]_net_1\, \RDATA_M_int_2[30]\, 
        \RDATA_M_int[31]_net_1\, \RDATA_M_int_2[31]\, 
        \RDATA_M_int[32]_net_1\, \RDATA_M_int_2[32]\, 
        \RDATA_M_int[3]_net_1\, \RDATA_M_int_2[3]\, 
        \RDATA_M_int[4]_net_1\, \RDATA_M_int_2[4]\, 
        \RDATA_M_int[5]_net_1\, \RDATA_M_int_2[5]\, 
        \RDATA_M_int[6]_net_1\, \RDATA_M_int_2[6]\, 
        \RDATA_M_int[7]_net_1\, \RDATA_M_int_2[7]\, 
        \RDATA_M_int[8]_net_1\, \RDATA_M_int_2[8]\, 
        \RDATA_M_int[9]_net_1\, \RDATA_M_int_2[9]\, 
        \RDATA_M_int[10]_net_1\, \RDATA_M_int_2[10]\, 
        \RDATA_M_int[11]_net_1\, \RDATA_M_int_2[11]\, 
        \RDATA_M_int[12]_net_1\, \RDATA_M_int_2[12]\, 
        \RDATA_M_int[13]_net_1\, \RDATA_M_int_2[13]\, 
        \RDATA_M_int[14]_net_1\, \RDATA_M_int_2[14]\, 
        \RDATA_M_int[15]_net_1\, \RDATA_M_int_2[15]\, 
        \RDATA_M_int[16]_net_1\, \RDATA_M_int_2[16]\, 
        \RDATA_M_int[17]_net_1\, \RDATA_M_int_2[17]\, 
        \RDATA_M_int[0]_net_1\, \RDATA_M_int_2[0]\, 
        \RDATA_M_int[1]_net_1\, \RDATA_M_int_2[1]\, 
        \RDATA_M_int[2]_net_1\, \RDATA_M_int_2[2]\, 
        \WDATA_M_INPFF1[63]_net_1\, \wready_m_xhdl2\, 
        \WSTRB_M_INPFF1[0]_net_1\, \WSTRB_M_INPFF1[1]_net_1\, 
        \WSTRB_M_INPFF1[2]_net_1\, \WSTRB_M_INPFF1[3]_net_1\, 
        \WSTRB_M_INPFF1[4]_net_1\, \WSTRB_M_INPFF1[5]_net_1\, 
        \WSTRB_M_INPFF1[6]_net_1\, \WSTRB_M_INPFF1[7]_net_1\, 
        \WDATA_M_INPFF1[48]_net_1\, \WDATA_M_INPFF1[49]_net_1\, 
        \WDATA_M_INPFF1[50]_net_1\, \WDATA_M_INPFF1[51]_net_1\, 
        \WDATA_M_INPFF1[52]_net_1\, \WDATA_M_INPFF1[53]_net_1\, 
        \WDATA_M_INPFF1[54]_net_1\, \WDATA_M_INPFF1[55]_net_1\, 
        \WDATA_M_INPFF1[56]_net_1\, \WDATA_M_INPFF1[57]_net_1\, 
        \WDATA_M_INPFF1[58]_net_1\, \WDATA_M_INPFF1[59]_net_1\, 
        \WDATA_M_INPFF1[60]_net_1\, \WDATA_M_INPFF1[61]_net_1\, 
        \WDATA_M_INPFF1[62]_net_1\, \WDATA_M_INPFF1[33]_net_1\, 
        \WDATA_M_INPFF1[34]_net_1\, \WDATA_M_INPFF1[35]_net_1\, 
        \WDATA_M_INPFF1[36]_net_1\, \WDATA_M_INPFF1[37]_net_1\, 
        \WDATA_M_INPFF1[38]_net_1\, \WDATA_M_INPFF1[39]_net_1\, 
        \WDATA_M_INPFF1[40]_net_1\, \WDATA_M_INPFF1[41]_net_1\, 
        \WDATA_M_INPFF1[42]_net_1\, \WDATA_M_INPFF1[43]_net_1\, 
        \WDATA_M_INPFF1[44]_net_1\, \WDATA_M_INPFF1[45]_net_1\, 
        \WDATA_M_INPFF1[46]_net_1\, \WDATA_M_INPFF1[47]_net_1\, 
        \WDATA_M_INPFF1[18]_net_1\, \WDATA_M_INPFF1[19]_net_1\, 
        \WDATA_M_INPFF1[20]_net_1\, \WDATA_M_INPFF1[21]_net_1\, 
        \WDATA_M_INPFF1[22]_net_1\, \WDATA_M_INPFF1[23]_net_1\, 
        \WDATA_M_INPFF1[24]_net_1\, \WDATA_M_INPFF1[25]_net_1\, 
        \WDATA_M_INPFF1[26]_net_1\, \WDATA_M_INPFF1[27]_net_1\, 
        \WDATA_M_INPFF1[28]_net_1\, \WDATA_M_INPFF1[29]_net_1\, 
        \WDATA_M_INPFF1[30]_net_1\, \WDATA_M_INPFF1[31]_net_1\, 
        \WDATA_M_INPFF1[32]_net_1\, \WDATA_M_INPFF1[3]_net_1\, 
        \WDATA_M_INPFF1[4]_net_1\, \WDATA_M_INPFF1[5]_net_1\, 
        \WDATA_M_INPFF1[6]_net_1\, \WDATA_M_INPFF1[7]_net_1\, 
        \WDATA_M_INPFF1[8]_net_1\, \WDATA_M_INPFF1[9]_net_1\, 
        \WDATA_M_INPFF1[10]_net_1\, \WDATA_M_INPFF1[11]_net_1\, 
        \WDATA_M_INPFF1[12]_net_1\, \WDATA_M_INPFF1[13]_net_1\, 
        \WDATA_M_INPFF1[14]_net_1\, \WDATA_M_INPFF1[15]_net_1\, 
        \WDATA_M_INPFF1[16]_net_1\, \WDATA_M_INPFF1[17]_net_1\, 
        \WDATA_M_INPFF1[0]_net_1\, \WDATA_M_INPFF1[1]_net_1\, 
        \WDATA_M_INPFF1[2]_net_1\, un2_arvalid_m, un2_awvalid_m, 
        \AWSIZE_M_INPFF1_3[0]\, \AWSIZE_M_INPFF1_3[1]\, 
        \ARSIZE_M_INPFF1_2[0]\, \ARSIZE_M_INPFF1_2[1]\, 
        \AWBURST_MI0[0]\, \prev_ARADDR[24]_net_1\, N_28_i, 
        \prev_ARADDR[25]_net_1\, \prev_ARADDR[26]_net_1\, 
        \prev_ARADDR[27]_net_1\, \rdtrans_inprog\, N_53, N_24, 
        \ARVALID_MI0\, N_28, \ARVALID_M_pulse_1_sqmuxa_i\, 
        \ARVALID_M_INPFF1\, N_12_i_0, \RVALID_M_int\, 
        RVALID_M_int_2, \RLAST_M_int\, RLAST_M_int_2, 
        \BVALID_M_pulse\, \BVALID_M_pulse_1_sqmuxa_i\, 
        \WVALID_M_pulse\, \WVALID_M_pulse_1_sqmuxa_i\, 
        \AWVALID_MI0\, \AWVALID_M_pulse_1_sqmuxa_i\, \WVALID_MI0\, 
        \WVALID_MI_xhdl25_2\, \COREAHBLTOAXI_0_AXIMasterIF_RLAST\, 
        RLAST_M_xhdl10_4, \COREAHBLTOAXI_0_AXIMasterIF_RVALID\, 
        RVALID_M_xhdl11_5, BVALID_M_xhdl5_5, \BVALID_M_INPFF1\, 
        BVALID_M_INPFF1_2, \add_rdtran\, 
        \un21_rlast_m_xhdl10_0_a2\, \stall_trans\, 
        \un23_arvalid_m_0_a2\, \temp_xhdl44\, \ARVALID_M_FF1\, 
        N_14_i_0, AWREADY_M_xhdl1_2, 
        \COREAHBLTOAXI_0_AXIMasterIF_WREADY\, WREADY_M_xhdl2_2, 
        \un36_rvalid_m_xhdl11\, \AWVALID_M_FF1\, AWVALID_M_FF1_2, 
        \WVALID_M_INPFF1\, WVALID_M_INPFF1_2, \WVALID_M_FF1\, 
        \BVALID_M_FF1\, \BVALID_IM_r\, N_32, N_22_i_1, N_29, N_81, 
        \RREADY_MI0\, \un21_arvalid_m_NE_1\, 
        \un21_arvalid_m_NE_0\, N_35, \SUM_i_0_tz[0]\, N_34, N_37, 
        N_41, \SUM_i_0_0[0]\, N_36 : std_logic;

begin 

    RREADY_MI0 <= \RREADY_MI0\;
    COREAHBLTOAXI_0_AXIMasterIF_WREADY <= 
        \COREAHBLTOAXI_0_AXIMasterIF_WREADY\;
    COREAHBLTOAXI_0_AXIMasterIF_RVALID <= 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\;
    COREAHBLTOAXI_0_AXIMasterIF_RLAST <= 
        \COREAHBLTOAXI_0_AXIMasterIF_RLAST\;
    WVALID_MI0 <= \WVALID_MI0\;
    AWVALID_MI0 <= \AWVALID_MI0\;
    ARVALID_MI0 <= \ARVALID_MI0\;
    wready_m_xhdl2 <= \wready_m_xhdl2\;
    COREAHBLTOAXI_0_AXIMasterIF_ARREADY <= 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\;
    COREAHBLTOAXI_0_AXIMasterIF_AWREADY <= 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\;
    COREAHBLTOAXI_0_AXIMasterIF_BVALID <= 
        \COREAHBLTOAXI_0_AXIMasterIF_BVALID\;

    \RDATA_M_int[63]\ : SLE
      port map(D => \RDATA_M_int_2[63]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[63]_net_1\);
    
    \RDATA_M_int[37]\ : SLE
      port map(D => \RDATA_M_int_2[37]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[37]_net_1\);
    
    \ARADDR_M_INPFF1[22]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(22));
    
    un21_rlast_m_xhdl10_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => \un36_rvalid_m_xhdl11\, B => N_28, Y => 
        \un21_rlast_m_xhdl10_0_a2\);
    
    \L5.RDATA_M_int_2[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(27), Y => 
        \RDATA_M_int_2[27]\);
    
    AWREADY_M_xhdl1 : SLE
      port map(D => AWREADY_M_xhdl1_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\);
    
    \WDATA_M_INPFF1[6]\ : SLE
      port map(D => N_278_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[6]_net_1\);
    
    \L5.RDATA_M_int_2[46]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(46), Y => 
        \RDATA_M_int_2[46]\);
    
    \WSTRB_M_INPFF1[6]\ : SLE
      port map(D => N_1451_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[6]_net_1\);
    
    \un1_rd_wdcntr_1_1.N_20_i\ : CFG4
      generic map(INIT => x"A965")

      port map(A => \rd_wdcntr[2]_net_1\, B => 
        \rd_wdcntr[1]_net_1\, C => N_35, D => N_32, Y => N_20_i);
    
    \RDATA_M_int[4]\ : SLE
      port map(D => \RDATA_M_int_2[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[4]_net_1\);
    
    \WDATA_M_INPFF1[7]\ : SLE
      port map(D => N_381_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[7]_net_1\);
    
    \WDATA_M_INPFF1[31]\ : SLE
      port map(D => N_195_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[31]_net_1\);
    
    \RDATA_M_xhdl8[59]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[59]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59));
    
    \RDATA_M_int[27]\ : SLE
      port map(D => \RDATA_M_int_2[27]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[27]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[27]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[27]_net_1\, Y
         => \RDATA_M_xhdl8_3[27]\);
    
    \ARADDR_M_INPFF1[13]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(13));
    
    \WDATA_MI_xhdl22[27]\ : SLE
      port map(D => \WDATA_M_INPFF1[27]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(27));
    
    \WDATA_M_INPFF1[59]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(59), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[59]_net_1\);
    
    \RDATA_M_xhdl8[52]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[52]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52));
    
    un21_arvalid_m_NE_0 : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \prev_ARADDR[27]_net_1\, B => 
        \prev_ARADDR[26]_net_1\, C => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), D => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), Y => 
        \un21_arvalid_m_NE_0\);
    
    \L5.RDATA_M_xhdl8_3[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[6]_net_1\, Y
         => \RDATA_M_xhdl8_3[6]\);
    
    \L3.WREADY_M_xhdl2_2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \WVALID_MI0\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_WREADY\, C => WREADY_IM0, Y
         => WREADY_M_xhdl2_2);
    
    BVALID_IM_r : SLE
      port map(D => BVALID_IM0, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \BVALID_IM_r\);
    
    \rd_wdcntr_RNIEOM[3]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rd_wdcntr[1]_net_1\, B => 
        \rd_wdcntr[3]_net_1\, Y => N_81);
    
    \L5.RDATA_M_int_2[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(0), Y => 
        \RDATA_M_int_2[0]\);
    
    \WDATA_MI_xhdl22[46]\ : SLE
      port map(D => \WDATA_M_INPFF1[46]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(46));
    
    \RDATA_M_xhdl8[23]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[23]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23));
    
    \L5.RDATA_M_xhdl8_3[57]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[57]_net_1\, Y
         => \RDATA_M_xhdl8_3[57]\);
    
    \AWADDR_M_INPFF1[15]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(15));
    
    \RDATA_M_xhdl8[56]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[56]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56));
    
    \AWBURST_M_INPFF1[0]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_AWREADY_i, CLK
         => SDRCLK_c, EN => N_75_i, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWBURST_MI0[0]\);
    
    \L5.RDATA_M_xhdl8_3[42]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[42]_net_1\, Y
         => \RDATA_M_xhdl8_3[42]\);
    
    \L5.RDATA_M_int_2[22]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(22), Y => 
        \RDATA_M_int_2[22]\);
    
    \RDATA_M_xhdl8[55]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[55]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55));
    
    \WDATA_M_INPFF1[10]\ : SLE
      port map(D => N_276_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[10]_net_1\);
    
    \WDATA_MI_xhdl22[57]\ : SLE
      port map(D => \WDATA_M_INPFF1[57]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(57));
    
    \RDATA_M_xhdl8[49]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[49]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49));
    
    \RDATA_M_xhdl8[28]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[28]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28));
    
    \L5.RLAST_M_int_2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RLAST_IM0, Y => 
        RLAST_M_int_2);
    
    \ARADDR_M_INPFF1[9]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(9));
    
    \WDATA_M_INPFF1[9]\ : SLE
      port map(D => N_277_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[9]_net_1\);
    
    \L5.RDATA_M_int_2[21]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(21), Y => 
        \RDATA_M_int_2[21]\);
    
    \RDATA_M_xhdl8[42]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[42]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42));
    
    \L5.RDATA_M_xhdl8_3[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[26]_net_1\, Y
         => \RDATA_M_xhdl8_3[26]\);
    
    BVALID_M_xhdl5 : SLE
      port map(D => BVALID_M_xhdl5_5, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_BVALID\);
    
    \ARADDR_M_INPFF1[8]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(8));
    
    \rd_wdcntr[1]\ : SLE
      port map(D => N_22_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rd_wdcntr[1]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[56]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[56]_net_1\, Y
         => \RDATA_M_xhdl8_3[56]\);
    
    \L5.RDATA_M_int_2[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(13), Y => 
        \RDATA_M_int_2[13]\);
    
    \AWBURST_M_INPFF1_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\, Y => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY_i);
    
    \ARSIZE_M_INPFF1[1]\ : SLE
      port map(D => \ARSIZE_M_INPFF1_2[1]\, CLK => SDRCLK_c, EN
         => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => ARSIZE_MI0(1));
    
    \RDATA_M_xhdl8[13]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[13]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13));
    
    \L5.RDATA_M_int_2[37]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(37), Y => 
        \RDATA_M_int_2[37]\);
    
    AWVALID_M_FF1 : SLE
      port map(D => AWVALID_M_FF1_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWVALID_M_FF1\);
    
    \RDATA_M_xhdl8[46]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[46]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46));
    
    \L5.RDATA_M_xhdl8_3[39]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[39]_net_1\, Y
         => \RDATA_M_xhdl8_3[39]\);
    
    \AWSIZE_M_INPFF1[1]\ : SLE
      port map(D => \AWSIZE_M_INPFF1_3[1]\, CLK => SDRCLK_c, EN
         => N_75_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWSIZE_MI0(1));
    
    \un1_rd_wdcntr_1_1.SUM_i_o2[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_35, B => \rd_wdcntr[1]_net_1\, Y => N_37);
    
    \ARADDR_M_INPFF1[27]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(27));
    
    \RDATA_M_xhdl8[7]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7));
    
    \RDATA_M_xhdl8[45]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[45]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45));
    
    \L3.AWREADY_M_xhdl1_2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \AWVALID_MI0\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\, C => AWREADY_IM0, 
        Y => AWREADY_M_xhdl1_2);
    
    \ARSIZE_M_INPFF1[0]\ : SLE
      port map(D => \ARSIZE_M_INPFF1_2[0]\, CLK => SDRCLK_c, EN
         => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => ARSIZE_MI0(0));
    
    \RDATA_M_int[6]\ : SLE
      port map(D => \RDATA_M_int_2[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[6]_net_1\);
    
    \WDATA_M_INPFF1[27]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(27), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[27]_net_1\);
    
    \L5.RDATA_M_int_2[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(8), Y => 
        \RDATA_M_int_2[8]\);
    
    \AWSIZE_M_INPFF1[0]\ : SLE
      port map(D => \AWSIZE_M_INPFF1_3[0]\, CLK => SDRCLK_c, EN
         => N_75_i, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWSIZE_MI0(0));
    
    RVALID_M_xhdl11 : SLE
      port map(D => RVALID_M_xhdl11_5, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\);
    
    \RDATA_M_xhdl8[18]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[18]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18));
    
    \L5.RDATA_M_int_2[57]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(57), Y => 
        \RDATA_M_int_2[57]\);
    
    RVALID_M_int : SLE
      port map(D => RVALID_M_int_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RVALID_M_int\);
    
    mst_wr_end : SLE
      port map(D => \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => m0_wr_end);
    
    \RDATA_M_int[46]\ : SLE
      port map(D => \RDATA_M_int_2[46]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[46]_net_1\);
    
    \WDATA_MI_xhdl22[17]\ : SLE
      port map(D => \WDATA_M_INPFF1[17]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(17));
    
    RLAST_M_xhdl10 : SLE
      port map(D => RLAST_M_xhdl10_4, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_RLAST\);
    
    \WDATA_MI_xhdl22[45]\ : SLE
      port map(D => \WDATA_M_INPFF1[45]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(45));
    
    \L5.RDATA_M_int_2[43]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(43), Y => 
        \RDATA_M_int_2[43]\);
    
    \AWADDR_M_INPFF1[21]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(21));
    
    \AWADDR_M_INPFF1[26]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(26));
    
    \WSTRB_M_INPFF1[1]\ : SLE
      port map(D => N_1446_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[1]_net_1\);
    
    \WDATA_MI_xhdl22[37]\ : SLE
      port map(D => \WDATA_M_INPFF1[37]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(37));
    
    \RDATA_M_int[0]\ : SLE
      port map(D => \RDATA_M_int_2[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[0]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[22]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[22]_net_1\, Y
         => \RDATA_M_xhdl8_3[22]\);
    
    \L5.RDATA_M_int_2[32]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(32), Y => 
        \RDATA_M_int_2[32]\);
    
    \ARADDR_M_INPFF1[7]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(7));
    
    \WDATA_M_INPFF1[50]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(50), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[50]_net_1\);
    
    \AWADDR_M_INPFF1[14]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(14));
    
    AWVALID_M_pulse : SLE
      port map(D => N_48, CLK => SDRCLK_c, EN => 
        \AWVALID_M_pulse_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWVALID_MI0\);
    
    \L5.RDATA_M_int_2[31]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(31), Y => 
        \RDATA_M_int_2[31]\);
    
    \WDATA_M_INPFF1[8]\ : SLE
      port map(D => N_382_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[8]_net_1\);
    
    \WDATA_M_INPFF1[23]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(23), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[23]_net_1\);
    
    \RDATA_M_int[42]\ : SLE
      port map(D => \RDATA_M_int_2[42]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[42]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[52]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[52]_net_1\, Y
         => \RDATA_M_xhdl8_3[52]\);
    
    \AWADDR_M_INPFF1[9]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(9));
    
    \WDATA_M_INPFF1[48]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(48), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[48]_net_1\);
    
    \un1_rd_wdcntr_1_1.SUM_i_0_0[0]\ : CFG4
      generic map(INIT => x"C30E")

      port map(A => \SUM_i_0_tz[0]\, B => \un36_rvalid_m_xhdl11\, 
        C => \rd_wdcntr[0]_net_1\, D => N_28, Y => \SUM_i_0_0[0]\);
    
    \L5.RDATA_M_xhdl8_3[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[7]_net_1\, Y
         => \RDATA_M_xhdl8_3[7]\);
    
    \L5.RDATA_M_int_2[52]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(52), Y => 
        \RDATA_M_int_2[52]\);
    
    \WSTRB_MI_xhdl23[6]\ : SLE
      port map(D => \WSTRB_M_INPFF1[6]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(6));
    
    un21_arvalid_m_NE_1 : CFG4
      generic map(INIT => x"7BDE")

      port map(A => \prev_ARADDR[25]_net_1\, B => 
        \prev_ARADDR[24]_net_1\, C => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25), D => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24), Y => 
        \un21_arvalid_m_NE_1\);
    
    \WDATA_MI_xhdl22[23]\ : SLE
      port map(D => \WDATA_M_INPFF1[23]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(23));
    
    \AWADDR_M_INPFF1[8]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(8));
    
    \L5.RDATA_M_int_2[51]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(51), Y => 
        \RDATA_M_int_2[51]\);
    
    ARVALID_M_INPFF1_RNO : CFG2
      generic map(INIT => x"1")

      port map(A => N_41, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => N_12_i_0);
    
    \rd_wdcntr[0]\ : SLE
      port map(D => N_16_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rd_wdcntr[0]_net_1\);
    
    \RDATA_M_xhdl8[33]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[33]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33));
    
    \L1.AWSIZE_M_INPFF1_3[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0), B => 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\, Y => 
        \AWSIZE_M_INPFF1_3[0]\);
    
    \L5.RDATA_M_int_2[28]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(28), Y => 
        \RDATA_M_int_2[28]\);
    
    \RDATA_M_int[34]\ : SLE
      port map(D => \RDATA_M_int_2[34]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[34]_net_1\);
    
    \ARADDR_M_INPFF1[19]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(19));
    
    \RDATA_M_int[48]\ : SLE
      port map(D => \RDATA_M_int_2[48]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[48]_net_1\);
    
    \L5.RDATA_M_int_2[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(10), Y => 
        \RDATA_M_int_2[10]\);
    
    \RDATA_M_xhdl8[2]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \WDATA_M_INPFF1[15]\ : SLE
      port map(D => N_203_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[15]_net_1\);
    
    \WDATA_MI_xhdl22[53]\ : SLE
      port map(D => \WDATA_M_INPFF1[53]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(53));
    
    \RDATA_M_xhdl8[38]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[38]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38));
    
    \RDATA_M_int[24]\ : SLE
      port map(D => \RDATA_M_int_2[24]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[24]_net_1\);
    
    \L5.RVALID_M_int_2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RVALID_IM0, Y => 
        RVALID_M_int_2);
    
    \WDATA_M_INPFF1[38]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(38), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[38]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[14]_net_1\, Y
         => \RDATA_M_xhdl8_3[14]\);
    
    \WDATA_MI_xhdl22[6]\ : SLE
      port map(D => \WDATA_M_INPFF1[6]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(6));
    
    \WDATA_MI_xhdl22[22]\ : SLE
      port map(D => \WDATA_M_INPFF1[22]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(22));
    
    stall_trans : SLE
      port map(D => \un23_arvalid_m_0_a2\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \stall_trans\);
    
    \RDATA_M_int[17]\ : SLE
      port map(D => \RDATA_M_int_2[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[17]_net_1\);
    
    ARREADY_M_xhdl6_RNI6A9T : CFG2
      generic map(INIT => x"8")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => N_28_i);
    
    \WDATA_MI_xhdl22[0]\ : SLE
      port map(D => \WDATA_M_INPFF1[0]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(0));
    
    \L5.RDATA_M_xhdl8_3[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[3]_net_1\, Y
         => \RDATA_M_xhdl8_3[3]\);
    
    \L5.RDATA_M_int_2[40]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(40), Y => 
        \RDATA_M_int_2[40]\);
    
    \AWADDR_M_INPFF1[7]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(7));
    
    \RDATA_M_xhdl8[4]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4));
    
    \L5.RDATA_M_int_2[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(5), Y => 
        \RDATA_M_int_2[5]\);
    
    \WDATA_M_INPFF1[24]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(24), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[24]_net_1\);
    
    \WDATA_M_INPFF1[16]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(16), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[16]_net_1\);
    
    \WDATA_MI_xhdl22[21]\ : SLE
      port map(D => \WDATA_M_INPFF1[21]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(21));
    
    un36_rvalid_m_xhdl11 : CFG2
      generic map(INIT => x"8")

      port map(A => \RREADY_MI0\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_RLAST\, Y => 
        \un36_rvalid_m_xhdl11\);
    
    \RDATA_M_xhdl8[53]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[53]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53));
    
    \RDATA_M_xhdl8[24]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[24]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24));
    
    \AWADDR_M_INPFF1[19]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(19));
    
    \AWADDR_M_INPFF1[18]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(18));
    
    \WDATA_MI_xhdl22[52]\ : SLE
      port map(D => \WDATA_M_INPFF1[52]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(52));
    
    \ARADDR_M_INPFF1[20]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(20));
    
    \RDATA_M_int[49]\ : SLE
      port map(D => \RDATA_M_int_2[49]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[49]_net_1\);
    
    \WDATA_MI_xhdl22[47]\ : SLE
      port map(D => \WDATA_M_INPFF1[47]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(47));
    
    \WDATA_MI_xhdl22[13]\ : SLE
      port map(D => \WDATA_M_INPFF1[13]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(13));
    
    \RDATA_M_int[35]\ : SLE
      port map(D => \RDATA_M_int_2[35]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[35]_net_1\);
    
    \L5.RDATA_M_int_2[38]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(38), Y => 
        \RDATA_M_int_2[38]\);
    
    \WDATA_M_INPFF1[63]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(63), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[63]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[33]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[33]_net_1\, Y
         => \RDATA_M_xhdl8_3[33]\);
    
    \RDATA_M_xhdl8[58]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[58]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58));
    
    \WDATA_MI_xhdl22[33]\ : SLE
      port map(D => \WDATA_M_INPFF1[33]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(33));
    
    \un1_rd_wdcntr_1_1.SUM_i_0_tz[0]\ : CFG3
      generic map(INIT => x"D5")

      port map(A => N_29, B => \rd_wdcntr[2]_net_1\, C => N_81, Y
         => \SUM_i_0_tz[0]\);
    
    \RDATA_M_int[31]\ : SLE
      port map(D => \RDATA_M_int_2[31]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[31]_net_1\);
    
    mst_rd_end : SLE
      port map(D => \un36_rvalid_m_xhdl11\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m0_rd_end);
    
    \WSTRB_M_INPFF1[5]\ : SLE
      port map(D => N_1450_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[5]_net_1\);
    
    \WDATA_M_INPFF1[29]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(29), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[29]_net_1\);
    
    \WDATA_MI_xhdl22[9]\ : SLE
      port map(D => \WDATA_M_INPFF1[9]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(9));
    
    \WDATA_MI_xhdl22[51]\ : SLE
      port map(D => \WDATA_M_INPFF1[51]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(51));
    
    \RDATA_M_int[25]\ : SLE
      port map(D => \RDATA_M_int_2[25]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[25]_net_1\);
    
    \WDATA_M_INPFF1[55]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(55), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[55]_net_1\);
    
    \RDATA_M_int[40]\ : SLE
      port map(D => \RDATA_M_int_2[40]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[40]_net_1\);
    
    \L5.RDATA_M_int_2[58]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(58), Y => 
        \RDATA_M_int_2[58]\);
    
    \RDATA_M_xhdl8[43]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[43]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43));
    
    \WDATA_M_INPFF1[12]\ : SLE
      port map(D => N_274_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[12]_net_1\);
    
    \ARADDR_M_INPFF1[26]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(26));
    
    \RDATA_M_int[21]\ : SLE
      port map(D => \RDATA_M_int_2[21]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[21]_net_1\);
    
    WVALID_MI_xhdl25 : SLE
      port map(D => \WVALID_MI_xhdl25_2\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WVALID_MI0\);
    
    \L5.RDATA_M_xhdl8_3[19]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[19]_net_1\, Y
         => \RDATA_M_xhdl8_3[19]\);
    
    \WDATA_MI_xhdl22[3]\ : SLE
      port map(D => \WDATA_M_INPFF1[3]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(3));
    
    \RDATA_M_xhdl8[14]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[14]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14));
    
    \WSTRB_MI_xhdl23[1]\ : SLE
      port map(D => \WSTRB_M_INPFF1[1]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(1));
    
    \rd_wdcntr[2]\ : SLE
      port map(D => N_20_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rd_wdcntr[2]_net_1\);
    
    \WDATA_M_INPFF1[0]\ : SLE
      port map(D => N_137_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[0]_net_1\);
    
    WVALID_M_INPFF1 : SLE
      port map(D => WVALID_M_INPFF1_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WVALID_M_INPFF1\);
    
    \RDATA_M_xhdl8[48]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[48]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48));
    
    \ARADDR_M_INPFF1[5]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(5));
    
    \L5.RDATA_M_int_2[19]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(19), Y => 
        \RDATA_M_int_2[19]\);
    
    \WDATA_M_INPFF1[47]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(47), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[47]_net_1\);
    
    \WDATA_MI_xhdl22[12]\ : SLE
      port map(D => \WDATA_M_INPFF1[12]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(12));
    
    \RDATA_M_int[57]\ : SLE
      port map(D => \RDATA_M_int_2[57]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[57]_net_1\);
    
    \RDATA_M_xhdl8[1]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1));
    
    \L5.RDATA_M_xhdl8_3[44]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[44]_net_1\, Y
         => \RDATA_M_xhdl8_3[44]\);
    
    \L5.RDATA_M_int_2[14]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(14), Y => 
        \RDATA_M_int_2[14]\);
    
    \WDATA_M_INPFF1[56]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(56), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[56]_net_1\);
    
    \WDATA_MI_xhdl22[32]\ : SLE
      port map(D => \WDATA_M_INPFF1[32]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(32));
    
    BVALID_M_FF1 : SLE
      port map(D => \BVALID_M_INPFF1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \BVALID_M_FF1\);
    
    \L5.RDATA_M_int_2[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(26), Y => 
        \RDATA_M_int_2[26]\);
    
    \AWADDR_M_INPFF1[12]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(12));
    
    \L5.RDATA_M_int_2[62]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(62), Y => 
        \RDATA_M_int_2[62]\);
    
    \WDATA_MI_xhdl22[11]\ : SLE
      port map(D => \WDATA_M_INPFF1[11]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(11));
    
    \un1_rd_wdcntr_1_1.SUM_i_o2[1]\ : CFG3
      generic map(INIT => x"DF")

      port map(A => \un36_rvalid_m_xhdl11\, B => 
        \rd_wdcntr[0]_net_1\, C => N_28, Y => N_35);
    
    \L5.RDATA_M_int_2[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(7), Y => 
        \RDATA_M_int_2[7]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \L5.RDATA_M_xhdl8_3[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[8]_net_1\, Y
         => \RDATA_M_xhdl8_3[8]\);
    
    \L5.RDATA_M_int_2[61]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(61), Y => 
        \RDATA_M_int_2[61]\);
    
    \WDATA_MI_xhdl22[31]\ : SLE
      port map(D => \WDATA_M_INPFF1[31]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(31));
    
    \WDATA_MI_xhdl22[60]\ : SLE
      port map(D => \WDATA_M_INPFF1[60]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(60));
    
    \RDATA_M_xhdl8[61]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[61]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61));
    
    \L5.RDATA_M_int_2[49]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(49), Y => 
        \RDATA_M_int_2[49]\);
    
    \WDATA_M_INPFF1[37]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(37), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[37]_net_1\);
    
    \L5.RDATA_M_int_2[44]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(44), Y => 
        \RDATA_M_int_2[44]\);
    
    \WDATA_M_INPFF1[43]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(43), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[43]_net_1\);
    
    \RDATA_M_xhdl8[60]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[60]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60));
    
    \WDATA_M_INPFF1[52]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(52), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[52]_net_1\);
    
    \RDATA_M_int[43]\ : SLE
      port map(D => \RDATA_M_int_2[43]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[43]_net_1\);
    
    \L5.RDATA_M_int_2[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(2), Y => 
        \RDATA_M_int_2[2]\);
    
    \rd_wdcntr_RNIQ2MA[2]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \rd_wdcntr[2]_net_1\, B => 
        \rd_wdcntr[0]_net_1\, C => N_81, D => 
        \un36_rvalid_m_xhdl11\, Y => N_53);
    
    ARVALID_M_pulse_1_sqmuxa_i : CFG4
      generic map(INIT => x"0F4F")

      port map(A => \ARVALID_M_FF1\, B => \ARVALID_M_INPFF1\, C
         => N_28, D => N_41, Y => \ARVALID_M_pulse_1_sqmuxa_i\);
    
    \un1_rd_wdcntr_1_1.N_22_i_1\ : CFG4
      generic map(INIT => x"2420")

      port map(A => N_28, B => \rd_wdcntr[0]_net_1\, C => 
        \un36_rvalid_m_xhdl11\, D => N_29, Y => N_22_i_1);
    
    \L5.RDATA_M_xhdl8_3[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[9]_net_1\, Y
         => \RDATA_M_xhdl8_3[9]\);
    
    \AWADDR_M_INPFF1[20]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(20));
    
    \un1_rd_wdcntr_1_1.SUM_i_o4[1]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_32, B => \rd_wdcntr[1]_net_1\, Y => N_36);
    
    \L5.RDATA_M_xhdl8_3[35]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[35]_net_1\, Y
         => \RDATA_M_xhdl8_3[35]\);
    
    \RDATA_M_xhdl8[34]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[34]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34));
    
    \RDATA_M_int[3]\ : SLE
      port map(D => \RDATA_M_int_2[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[3]_net_1\);
    
    \WDATA_M_INPFF1[20]\ : SLE
      port map(D => N_201_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[20]_net_1\);
    
    \RDATA_M_int[2]\ : SLE
      port map(D => \RDATA_M_int_2[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[2]_net_1\);
    
    \WDATA_M_INPFF1[11]\ : SLE
      port map(D => N_275_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[11]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[30]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[30]_net_1\, Y
         => \RDATA_M_xhdl8_3[30]\);
    
    \WSTRB_M_INPFF1[4]\ : SLE
      port map(D => N_1449_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[4]_net_1\);
    
    \WDATA_MI_xhdl22[43]\ : SLE
      port map(D => \WDATA_M_INPFF1[43]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(43));
    
    \RDATA_M_int[36]\ : SLE
      port map(D => \RDATA_M_int_2[36]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[36]_net_1\);
    
    \RDATA_M_int[14]\ : SLE
      port map(D => \RDATA_M_int_2[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[14]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[24]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[24]_net_1\, Y
         => \RDATA_M_xhdl8_3[24]\);
    
    \AWADDR_M_INPFF1[5]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(5));
    
    \AWADDR_M_INPFF1[23]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(23));
    
    \WDATA_M_INPFF1[33]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(33), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[33]_net_1\);
    
    \RDATA_M_xhdl8[21]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[21]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21));
    
    ARVALID_M_pulse : SLE
      port map(D => N_28, CLK => SDRCLK_c, EN => 
        \ARVALID_M_pulse_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ARVALID_MI0\);
    
    \ARADDR_M_INPFF1[12]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(12));
    
    \L5.RDATA_M_int_2[36]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(36), Y => 
        \RDATA_M_int_2[36]\);
    
    BVALID_M_INPFF1 : SLE
      port map(D => BVALID_M_INPFF1_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \BVALID_M_INPFF1\);
    
    \WDATA_MI_xhdl22[24]\ : SLE
      port map(D => \WDATA_M_INPFF1[24]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(24));
    
    \L5.RDATA_M_xhdl8_3[49]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[49]_net_1\, Y
         => \RDATA_M_xhdl8_3[49]\);
    
    \RDATA_M_int[26]\ : SLE
      port map(D => \RDATA_M_int_2[26]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[26]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[54]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[54]_net_1\, Y
         => \RDATA_M_xhdl8_3[54]\);
    
    \ARADDR_M_INPFF1[4]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(4));
    
    \RDATA_M_xhdl8[20]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[20]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20));
    
    \L1.wready_m_xhdl2\ : CFG2
      generic map(INIT => x"7")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_WREADY\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, Y => \wready_m_xhdl2\);
    
    \WSTRB_M_INPFF1[3]\ : SLE
      port map(D => N_1448_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[3]_net_1\);
    
    \RDATA_M_int[32]\ : SLE
      port map(D => \RDATA_M_int_2[32]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[32]_net_1\);
    
    \L5.RDATA_M_int_2[56]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(56), Y => 
        \RDATA_M_int_2[56]\);
    
    RREADY_MI : CFG2
      generic map(INIT => x"8")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_RREADY, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\, Y => \RREADY_MI0\);
    
    \ARADDR_M_INPFF1[21]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(21));
    
    \L5.RDATA_M_xhdl8_3[63]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[63]_net_1\, Y
         => \RDATA_M_xhdl8_3[63]\);
    
    \L5.RDATA_M_int_2[23]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(23), Y => 
        \RDATA_M_int_2[23]\);
    
    ARVALID_M_INPFF1 : SLE
      port map(D => N_12_i_0, CLK => SDRCLK_c, EN => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \ARVALID_M_INPFF1\);
    
    \WDATA_M_INPFF1[44]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(44), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[44]_net_1\);
    
    \WDATA_MI_xhdl22[54]\ : SLE
      port map(D => \WDATA_M_INPFF1[54]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(54));
    
    \RDATA_M_int[22]\ : SLE
      port map(D => \RDATA_M_int_2[22]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[22]_net_1\);
    
    \WDATA_MI_xhdl22[42]\ : SLE
      port map(D => \WDATA_M_INPFF1[42]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(42));
    
    \RDATA_M_xhdl8[54]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[54]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54));
    
    \RDATA_M_xhdl8[11]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[11]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11));
    
    \RDATA_M_int[38]\ : SLE
      port map(D => \RDATA_M_int_2[38]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[38]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[13]_net_1\, Y
         => \RDATA_M_xhdl8_3[13]\);
    
    \L1.un2_awvalid_m\ : CFG3
      generic map(INIT => x"08")

      port map(A => axi_current_state_3, B => N_48, C => 
        awaddr_awvalid_clr_d, Y => un2_awvalid_m);
    
    \RDATA_M_xhdl8[10]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[10]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10));
    
    \L5.RDATA_M_xhdl8_3[31]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[31]_net_1\, Y
         => \RDATA_M_xhdl8_3[31]\);
    
    \WDATA_M_INPFF1[51]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(51), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[51]_net_1\);
    
    \WDATA_MI_xhdl22[41]\ : SLE
      port map(D => \WDATA_M_INPFF1[41]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(41));
    
    \RDATA_M_int[15]\ : SLE
      port map(D => \RDATA_M_int_2[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[15]_net_1\);
    
    \L5.RDATA_M_int_2[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(15), Y => 
        \RDATA_M_int_2[15]\);
    
    \RDATA_M_int[28]\ : SLE
      port map(D => \RDATA_M_int_2[28]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[28]_net_1\);
    
    \ARLOCK_M_INPFF1[1]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, CLK => 
        SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ARLOCK_MI0[1]\);
    
    \un1_rd_wdcntr_1_1.SUM_i_o2[0]\ : CFG3
      generic map(INIT => x"37")

      port map(A => \un21_arvalid_m_NE_0\, B => \rdtrans_inprog\, 
        C => \un21_arvalid_m_NE_1\, Y => N_29);
    
    \L5.BVALID_M_xhdl5_5\ : CFG2
      generic map(INIT => x"4")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, B => 
        \BVALID_M_pulse\, Y => BVALID_M_xhdl5_5);
    
    \WDATA_M_INPFF1[49]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(49), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[49]_net_1\);
    
    \AWADDR_M_INPFF1[27]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(27));
    
    \WDATA_M_INPFF1[34]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(34), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[34]_net_1\);
    
    \RDATA_M_int[54]\ : SLE
      port map(D => \RDATA_M_int_2[54]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[54]_net_1\);
    
    \RDATA_M_int[11]\ : SLE
      port map(D => \RDATA_M_int_2[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[11]_net_1\);
    
    \RDATA_M_xhdl8[8]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8));
    
    \L5.RDATA_M_xhdl8_3[29]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[29]_net_1\, Y
         => \RDATA_M_xhdl8_3[29]\);
    
    un23_arvalid_m_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => N_29, B => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, Y => 
        \un23_arvalid_m_0_a2\);
    
    \un1_rd_wdcntr_1_1.N_22_i\ : CFG4
      generic map(INIT => x"73C0")

      port map(A => N_28, B => \rd_wdcntr[1]_net_1\, C => N_32, D
         => N_22_i_1, Y => N_22_i);
    
    \RDATA_M_xhdl8[44]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[44]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44));
    
    \WDATA_M_INPFF1[60]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(60), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[60]_net_1\);
    
    \ARADDR_M_INPFF1[17]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(17));
    
    \L5.RDATA_M_xhdl8_3[38]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[38]_net_1\, Y
         => \RDATA_M_xhdl8_3[38]\);
    
    \WDATA_MI_xhdl22[4]\ : SLE
      port map(D => \WDATA_M_INPFF1[4]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(4));
    
    \AWADDR_M_INPFF1[4]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(4));
    
    \WDATA_MI_xhdl22[14]\ : SLE
      port map(D => \WDATA_M_INPFF1[14]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(14));
    
    \L5.RDATA_M_xhdl8_3[59]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[59]_net_1\, Y
         => \RDATA_M_xhdl8_3[59]\);
    
    \WSTRB_MI_xhdl23[4]\ : SLE
      port map(D => \WSTRB_M_INPFF1[4]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(4));
    
    \WDATA_MI_xhdl22[34]\ : SLE
      port map(D => \WDATA_M_INPFF1[34]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(34));
    
    \L5.RDATA_M_int_2[45]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(45), Y => 
        \RDATA_M_int_2[45]\);
    
    \RDATA_M_xhdl8[3]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3));
    
    \ARADDR_M_INPFF1[14]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(14));
    
    \WDATA_M_INPFF1[2]\ : SLE
      port map(D => N_135_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[2]_net_1\);
    
    \L5.RDATA_M_int_2[33]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(33), Y => 
        \RDATA_M_int_2[33]\);
    
    \WDATA_M_INPFF1[25]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(25), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[25]_net_1\);
    
    \WDATA_M_INPFF1[39]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(39), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[39]_net_1\);
    
    \AWADDR_M_INPFF1[11]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(11));
    
    \ARADDR_M_INPFF1[6]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(6));
    
    \AWADDR_M_INPFF1[16]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(16));
    
    \RDATA_M_int[39]\ : SLE
      port map(D => \RDATA_M_int_2[39]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[39]_net_1\);
    
    \WDATA_M_INPFF1[5]\ : SLE
      port map(D => N_380_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[5]_net_1\);
    
    \RDATA_M_xhdl8[31]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[31]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31));
    
    \L5.RDATA_M_int_2[20]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(20), Y => 
        \RDATA_M_int_2[20]\);
    
    \L5.RDATA_M_int_2[53]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(53), Y => 
        \RDATA_M_int_2[53]\);
    
    \ARBURST_M_INPFF1_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY_i);
    
    \RDATA_M_int[29]\ : SLE
      port map(D => \RDATA_M_int_2[29]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[29]_net_1\);
    
    \L1.WVALID_M_INPFF1_2\ : CFG2
      generic map(INIT => x"4")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_WREADY\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, Y => 
        WVALID_M_INPFF1_2);
    
    \RDATA_M_int[30]\ : SLE
      port map(D => \RDATA_M_int_2[30]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[30]_net_1\);
    
    temp_xhdl44 : CFG4
      generic map(INIT => x"1000")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, B => 
        N_41, C => ARREADY_IM0, D => \ARVALID_MI0\, Y => 
        \temp_xhdl44\);
    
    \RDATA_M_xhdl8[30]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[30]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30));
    
    \RDATA_M_xhdl8[0]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0));
    
    \L5.RDATA_M_xhdl8_3[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[2]_net_1\, Y
         => \RDATA_M_xhdl8_3[2]\);
    
    \L1.AWSIZE_M_INPFF1_3[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1), B => 
        \COREAHBLTOAXI_0_AXIMasterIF_AWREADY\, Y => 
        \AWSIZE_M_INPFF1_3[1]\);
    
    \WDATA_M_INPFF1[26]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(26), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[26]_net_1\);
    
    \RDATA_M_int[55]\ : SLE
      port map(D => \RDATA_M_int_2[55]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[55]_net_1\);
    
    \WDATA_M_INPFF1[18]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(18), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[18]_net_1\);
    
    \RDATA_M_xhdl8[5]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5));
    
    \RDATA_M_int[20]\ : SLE
      port map(D => \RDATA_M_int_2[20]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[20]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[60]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[60]_net_1\, Y
         => \RDATA_M_xhdl8_3[60]\);
    
    \L5.RDATA_M_xhdl8_3[37]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[37]_net_1\, Y
         => \RDATA_M_xhdl8_3[37]\);
    
    \ARADDR_M_INPFF1[23]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(23));
    
    \WDATA_MI_xhdl22[28]\ : SLE
      port map(D => \WDATA_M_INPFF1[28]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(28));
    
    \AWLOCK_M_INPFF1_RNIFGIE[1]\ : CFG1
      generic map(INIT => "01")

      port map(A => \AWLOCK_MI0[1]\, Y => AWLOCK_MI0_i_0);
    
    \RDATA_M_int[51]\ : SLE
      port map(D => \RDATA_M_int_2[51]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[51]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[43]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[43]_net_1\, Y
         => \RDATA_M_xhdl8_3[43]\);
    
    \L1.un2_arvalid_m_0_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => un2_arvalid_m);
    
    \RDATA_M_int[61]\ : SLE
      port map(D => \RDATA_M_int_2[61]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[61]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[15]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[15]_net_1\, Y
         => \RDATA_M_xhdl8_3[15]\);
    
    \WDATA_M_INPFF1[40]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(40), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[40]_net_1\);
    
    \ARADDR_M_INPFF1[15]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(15));
    
    \WSTRB_M_INPFF1[7]\ : SLE
      port map(D => N_1452_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[7]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[10]_net_1\, Y
         => \RDATA_M_xhdl8_3[10]\);
    
    BVALID_M_pulse : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_BVALID_i, CLK => 
        SDRCLK_c, EN => \BVALID_M_pulse_1_sqmuxa_i\, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \BVALID_M_pulse\);
    
    AWVALID_M_pulse_1_sqmuxa_i : CFG3
      generic map(INIT => x"4F")

      port map(A => \AWVALID_M_FF1\, B => \AWBURST_MI0[0]\, C => 
        N_48, Y => \AWVALID_M_pulse_1_sqmuxa_i\);
    
    RLAST_M_int : SLE
      port map(D => RLAST_M_int_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RLAST_M_int\);
    
    \L5.RDATA_M_int_2[17]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(17), Y => 
        \RDATA_M_int_2[17]\);
    
    rdtrans_inprog_1_sqmuxa_i_0 : CFG3
      generic map(INIT => x"BF")

      port map(A => \add_rdtran\, B => N_28, C => N_53, Y => N_24);
    
    \WSTRB_M_INPFF1[2]\ : SLE
      port map(D => N_1447_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[2]_net_1\);
    
    \WSTRB_MI_xhdl23[0]\ : SLE
      port map(D => \WSTRB_M_INPFF1[0]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(0));
    
    \WDATA_MI_xhdl22[58]\ : SLE
      port map(D => \WDATA_M_INPFF1[58]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(58));
    
    \RDATA_M_xhdl8[51]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[51]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51));
    
    \RDATA_M_int[16]\ : SLE
      port map(D => \RDATA_M_int_2[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[16]_net_1\);
    
    \WDATA_M_INPFF1[22]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(22), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[22]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[36]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[36]_net_1\, Y
         => \RDATA_M_xhdl8_3[36]\);
    
    \AWADDR_M_INPFF1[6]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(6));
    
    \un1_rd_wdcntr_1_1.SUM_i_o4[0]\ : CFG4
      generic map(INIT => x"FBFF")

      port map(A => N_28, B => \rd_wdcntr[0]_net_1\, C => 
        \un36_rvalid_m_xhdl11\, D => N_29, Y => N_32);
    
    \L5.RDATA_M_int_2[30]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(30), Y => 
        \RDATA_M_int_2[30]\);
    
    \L1.ARVALID_M_FF1_2_i_o2\ : CFG4
      generic map(INIT => x"20FF")

      port map(A => \rd_wdcntr[2]_net_1\, B => 
        \rd_wdcntr[0]_net_1\, C => N_81, D => N_29, Y => N_34);
    
    \RDATA_M_xhdl8[50]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[50]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50));
    
    \RDATA_M_xhdl8[27]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[27]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27));
    
    \WSTRB_MI_xhdl23[5]\ : SLE
      port map(D => \WSTRB_M_INPFF1[5]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(5));
    
    \RDATA_M_xhdl8[6]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6));
    
    \RDATA_M_int[8]\ : SLE
      port map(D => \RDATA_M_int_2[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[8]_net_1\);
    
    \ARBURST_M_INPFF1[0]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARREADY_i, CLK
         => SDRCLK_c, EN => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => ARBURST_MI0_0);
    
    \ARLOCK_M_INPFF1_RNIA0OB[1]\ : CFG1
      generic map(INIT => "01")

      port map(A => \ARLOCK_MI0[1]\, Y => ARLOCK_MI0_i_0);
    
    \WDATA_M_INPFF1[30]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(30), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[30]_net_1\);
    
    \RDATA_M_int[1]\ : SLE
      port map(D => \RDATA_M_int_2[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[1]_net_1\);
    
    \ARADDR_M_INPFF1[3]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(3));
    
    \WDATA_MI_xhdl22[44]\ : SLE
      port map(D => \WDATA_M_INPFF1[44]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(44));
    
    \WDATA_MI_xhdl22[1]\ : SLE
      port map(D => \WDATA_M_INPFF1[1]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(1));
    
    \RDATA_M_int[33]\ : SLE
      port map(D => \RDATA_M_int_2[33]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[33]_net_1\);
    
    \L5.RDATA_M_int_2[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(4), Y => 
        \RDATA_M_int_2[4]\);
    
    \L5.RDATA_M_int_2[47]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(47), Y => 
        \RDATA_M_int_2[47]\);
    
    \RDATA_M_int[12]\ : SLE
      port map(D => \RDATA_M_int_2[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[12]_net_1\);
    
    \L5.RDATA_M_int_2[50]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(50), Y => 
        \RDATA_M_int_2[50]\);
    
    ARVALID_M_FF1 : SLE
      port map(D => N_14_i_0, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ARVALID_M_FF1\);
    
    add_rdtran : SLE
      port map(D => \un21_rlast_m_xhdl10_0_a2\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \add_rdtran\);
    
    \RDATA_M_xhdl8[41]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[41]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41));
    
    \L5.RDATA_M_xhdl8_3[61]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[61]_net_1\, Y
         => \RDATA_M_xhdl8_3[61]\);
    
    \L5.RDATA_M_int_2[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(12), Y => 
        \RDATA_M_int_2[12]\);
    
    \WDATA_M_INPFF1[58]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(58), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[58]_net_1\);
    
    \WDATA_MI_xhdl22[29]\ : SLE
      port map(D => \WDATA_M_INPFF1[29]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(29));
    
    \L5.RVALID_M_xhdl11_5\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RVALID_M_int\, Y => 
        RVALID_M_xhdl11_5);
    
    \ARADDR_M_INPFF1[10]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(10));
    
    \RDATA_M_int[23]\ : SLE
      port map(D => \RDATA_M_int_2[23]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[23]_net_1\);
    
    \L5.RDATA_M_int_2[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(11), Y => 
        \RDATA_M_int_2[11]\);
    
    \L5.RDATA_M_xhdl8_3[23]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[23]_net_1\, Y
         => \RDATA_M_xhdl8_3[23]\);
    
    \RDATA_M_xhdl8[40]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[40]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40));
    
    \L5.RDATA_M_int_2[29]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(29), Y => 
        \RDATA_M_int_2[29]\);
    
    WVALID_M_pulse : SLE
      port map(D => \wready_m_xhdl2\, CLK => SDRCLK_c, EN => 
        \WVALID_M_pulse_1_sqmuxa_i\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \WVALID_M_pulse\);
    
    \WDATA_MI_xhdl22[18]\ : SLE
      port map(D => \WDATA_M_INPFF1[18]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(18));
    
    \L5.RDATA_M_int_2[24]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(24), Y => 
        \RDATA_M_int_2[24]\);
    
    \RDATA_M_xhdl8[17]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[17]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17));
    
    \RDATA_M_int[18]\ : SLE
      port map(D => \RDATA_M_int_2[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[18]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[11]_net_1\, Y
         => \RDATA_M_xhdl8_3[11]\);
    
    \RDATA_M_int[47]\ : SLE
      port map(D => \RDATA_M_int_2[47]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[47]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[53]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[53]_net_1\, Y
         => \RDATA_M_xhdl8_3[53]\);
    
    WVALID_MI_xhdl25_2 : CFG2
      generic map(INIT => x"8")

      port map(A => \wready_m_xhdl2\, B => \WVALID_M_pulse\, Y
         => \WVALID_MI_xhdl25_2\);
    
    \WDATA_M_INPFF1[3]\ : SLE
      port map(D => N_134_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[3]_net_1\);
    
    \WDATA_MI_xhdl22[38]\ : SLE
      port map(D => \WDATA_M_INPFF1[38]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(38));
    
    \WDATA_MI_xhdl22[20]\ : SLE
      port map(D => \WDATA_M_INPFF1[20]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(20));
    
    \L5.RDATA_M_xhdl8_3[32]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[32]_net_1\, Y
         => \RDATA_M_xhdl8_3[32]\);
    
    \WDATA_MI_xhdl22[59]\ : SLE
      port map(D => \WDATA_M_INPFF1[59]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(59));
    
    \un1_rd_wdcntr_1_1.N_16_i\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_32, B => \SUM_i_0_0[0]\, Y => N_16_i);
    
    \ARADDR_M_INPFF1[16]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(16));
    
    \L5.RLAST_M_xhdl10_4\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RLAST_M_int\, Y => 
        RLAST_M_xhdl10_4);
    
    \L5.RDATA_M_int_2[42]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(42), Y => 
        \RDATA_M_int_2[42]\);
    
    \L5.RDATA_M_int_2[41]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(41), Y => 
        \RDATA_M_int_2[41]\);
    
    BVALID_M_pulse_1_sqmuxa_i : CFG3
      generic map(INIT => x"CE")

      port map(A => \BVALID_M_INPFF1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, C => \BVALID_M_FF1\, 
        Y => \BVALID_M_pulse_1_sqmuxa_i\);
    
    \RDATA_M_int[56]\ : SLE
      port map(D => \RDATA_M_int_2[56]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[56]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[45]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[45]_net_1\, Y
         => \RDATA_M_xhdl8_3[45]\);
    
    \L5.RDATA_M_xhdl8_3[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[18]_net_1\, Y
         => \RDATA_M_xhdl8_3[18]\);
    
    \L1.AWVALID_M_FF1_2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_48, B => \AWBURST_MI0[0]\, Y => 
        AWVALID_M_FF1_2);
    
    \L5.RDATA_M_xhdl8_3[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[1]_net_1\, Y
         => \RDATA_M_xhdl8_3[1]\);
    
    \rd_wdcntr[3]\ : SLE
      port map(D => N_18_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rd_wdcntr[3]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[40]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[40]_net_1\, Y
         => \RDATA_M_xhdl8_3[40]\);
    
    WVALID_M_FF1 : SLE
      port map(D => \WVALID_M_INPFF1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WVALID_M_FF1\);
    
    \RDATA_M_xhdl8[62]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[62]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62));
    
    \WDATA_M_INPFF1[62]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(62), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[62]_net_1\);
    
    \WDATA_M_INPFF1[21]\ : SLE
      port map(D => N_200_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[21]_net_1\);
    
    \WDATA_MI_xhdl22[50]\ : SLE
      port map(D => \WDATA_M_INPFF1[50]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(50));
    
    \L5.RDATA_M_int_2[63]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(63), Y => 
        \RDATA_M_int_2[63]\);
    
    \WDATA_M_INPFF1[17]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(17), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[17]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[5]_net_1\, Y
         => \RDATA_M_xhdl8_3[5]\);
    
    \L5.RDATA_M_int_2[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(9), Y => 
        \RDATA_M_int_2[9]\);
    
    \AWADDR_M_INPFF1[3]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(3));
    
    \WDATA_M_INPFF1[45]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(45), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[45]_net_1\);
    
    \RDATA_M_int[52]\ : SLE
      port map(D => \RDATA_M_int_2[52]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[52]_net_1\);
    
    \prev_ARADDR[25]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25), CLK
         => SDRCLK_c, EN => N_28_i, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \prev_ARADDR[25]_net_1\);
    
    \RDATA_M_int[62]\ : SLE
      port map(D => \RDATA_M_int_2[62]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[62]_net_1\);
    
    \RDATA_M_int[19]\ : SLE
      port map(D => \RDATA_M_int_2[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[19]_net_1\);
    
    \L5.RDATA_M_int_2[39]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(39), Y => 
        \RDATA_M_int_2[39]\);
    
    \WDATA_MI_xhdl22[19]\ : SLE
      port map(D => \WDATA_M_INPFF1[19]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(19));
    
    \WSTRB_MI_xhdl23[3]\ : SLE
      port map(D => \WSTRB_M_INPFF1[3]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(3));
    
    \L5.RDATA_M_int_2[34]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(34), Y => 
        \RDATA_M_int_2[34]\);
    
    ARVALID_M_FF1_RNO : CFG3
      generic map(INIT => x"08")

      port map(A => \ARVALID_M_INPFF1\, B => N_28, C => N_34, Y
         => N_14_i_0);
    
    \WDATA_MI_xhdl22[26]\ : SLE
      port map(D => \WDATA_M_INPFF1[26]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(26));
    
    \WDATA_MI_xhdl22[39]\ : SLE
      port map(D => \WDATA_M_INPFF1[39]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(39));
    
    \RDATA_M_int[9]\ : SLE
      port map(D => \RDATA_M_int_2[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[9]_net_1\);
    
    \RDATA_M_xhdl8[37]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[37]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37));
    
    \RDATA_M_xhdl8[29]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[29]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29));
    
    \RDATA_M_int[58]\ : SLE
      port map(D => \RDATA_M_int_2[58]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[58]_net_1\);
    
    \RDATA_M_int[10]\ : SLE
      port map(D => \RDATA_M_int_2[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[10]_net_1\);
    
    \L5.RDATA_M_int_2[59]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(59), Y => 
        \RDATA_M_int_2[59]\);
    
    \WDATA_M_INPFF1[46]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(46), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[46]_net_1\);
    
    \L5.RDATA_M_int_2[18]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(18), Y => 
        \RDATA_M_int_2[18]\);
    
    \RDATA_M_xhdl8[22]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[22]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22));
    
    \L5.RDATA_M_int_2[54]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(54), Y => 
        \RDATA_M_int_2[54]\);
    
    \WDATA_M_INPFF1[35]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(35), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[35]_net_1\);
    
    \WDATA_M_INPFF1[13]\ : SLE
      port map(D => N_273_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[13]_net_1\);
    
    \WDATA_MI_xhdl22[63]\ : SLE
      port map(D => \WDATA_M_INPFF1[63]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(63));
    
    \L5.RDATA_M_xhdl8_3[17]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[17]_net_1\, Y
         => \RDATA_M_xhdl8_3[17]\);
    
    \AWADDR_M_INPFF1[10]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(10));
    
    \WDATA_MI_xhdl22[10]\ : SLE
      port map(D => \WDATA_M_INPFF1[10]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(10));
    
    \L5.RDATA_M_xhdl8_3[25]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[25]_net_1\, Y
         => \RDATA_M_xhdl8_3[25]\);
    
    BVALID_M_pulse_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, Y => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID_i);
    
    \WDATA_MI_xhdl22[56]\ : SLE
      port map(D => \WDATA_M_INPFF1[56]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(56));
    
    \WDATA_MI_xhdl22[30]\ : SLE
      port map(D => \WDATA_M_INPFF1[30]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(30));
    
    \L5.RDATA_M_xhdl8_3[41]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[41]_net_1\, Y
         => \RDATA_M_xhdl8_3[41]\);
    
    \L5.RDATA_M_xhdl8_3[20]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[20]_net_1\, Y
         => \RDATA_M_xhdl8_3[20]\);
    
    \RDATA_M_xhdl8[26]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[26]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26));
    
    ARREADY_M_xhdl6_RNINF451 : CFG3
      generic map(INIT => x"BF")

      port map(A => araddr_arvalid_clr_d, B => 
        axi_current_state_0, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => N_28);
    
    \WDATA_MI_xhdl22[5]\ : SLE
      port map(D => \WDATA_M_INPFF1[5]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(5));
    
    \L5.RDATA_M_xhdl8_3[55]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[55]_net_1\, Y
         => \RDATA_M_xhdl8_3[55]\);
    
    \RDATA_M_xhdl8[25]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[25]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25));
    
    \AWADDR_M_INPFF1[13]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(13));
    
    ARREADY_M_xhdl6 : SLE
      port map(D => \temp_xhdl44\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\);
    
    \WDATA_M_INPFF1[57]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(57), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[57]_net_1\);
    
    \WDATA_MI_xhdl22[48]\ : SLE
      port map(D => \WDATA_M_INPFF1[48]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(48));
    
    \L5.RDATA_M_xhdl8_3[50]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[50]_net_1\, Y
         => \RDATA_M_xhdl8_3[50]\);
    
    \WREADY_M_xhdl2\ : SLE
      port map(D => WREADY_M_xhdl2_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_WREADY\);
    
    \L5.RDATA_M_int_2[48]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(48), Y => 
        \RDATA_M_int_2[48]\);
    
    \L1.BVALID_M_INPFF1_2\ : CFG3
      generic map(INIT => x"04")

      port map(A => \BVALID_IM_r\, B => BVALID_IM0, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_BVALID\, Y => 
        BVALID_M_INPFF1_2);
    
    \ARADDR_M_INPFF1[2]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(2));
    
    \WDATA_M_INPFF1[36]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(36), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[36]_net_1\);
    
    \RDATA_M_xhdl8[19]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[19]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19));
    
    \L1.ARSIZE_M_INPFF1_2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0), B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => 
        \ARSIZE_M_INPFF1_2[0]\);
    
    \WDATA_M_INPFF1[42]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(42), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[42]_net_1\);
    
    \prev_ARADDR[24]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24), CLK
         => SDRCLK_c, EN => N_28_i, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \prev_ARADDR[24]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[48]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[48]_net_1\, Y
         => \RDATA_M_xhdl8_3[48]\);
    
    \L5.RDATA_M_int_2[60]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(60), Y => 
        \RDATA_M_int_2[60]\);
    
    \WDATA_MI_xhdl22[7]\ : SLE
      port map(D => \WDATA_M_INPFF1[7]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(7));
    
    \RDATA_M_xhdl8[12]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[12]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12));
    
    \L5.RDATA_M_xhdl8_3[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[16]_net_1\, Y
         => \RDATA_M_xhdl8_3[16]\);
    
    \WDATA_M_INPFF1[61]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(61), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[61]_net_1\);
    
    \WDATA_MI_xhdl22[62]\ : SLE
      port map(D => \WDATA_M_INPFF1[62]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(62));
    
    \RDATA_M_xhdl8[57]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[57]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57));
    
    \L5.RDATA_M_int_2[25]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(25), Y => 
        \RDATA_M_int_2[25]\);
    
    \L5.RDATA_M_int_2[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(3), Y => 
        \RDATA_M_int_2[3]\);
    
    \ARADDR_M_INPFF1[11]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(11));
    
    \RDATA_M_int[59]\ : SLE
      port map(D => \RDATA_M_int_2[59]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[59]_net_1\);
    
    WVALID_M_pulse_1_sqmuxa_i : CFG3
      generic map(INIT => x"3B")

      port map(A => \WVALID_M_INPFF1\, B => \wready_m_xhdl2\, C
         => \WVALID_M_FF1\, Y => \WVALID_M_pulse_1_sqmuxa_i\);
    
    \WDATA_MI_xhdl22[25]\ : SLE
      port map(D => \WDATA_M_INPFF1[25]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(25));
    
    \RDATA_M_xhdl8[16]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[16]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16));
    
    \WDATA_MI_xhdl22[16]\ : SLE
      port map(D => \WDATA_M_INPFF1[16]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(16));
    
    \RDATA_M_xhdl8[15]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[15]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15));
    
    \WDATA_MI_xhdl22[61]\ : SLE
      port map(D => \WDATA_M_INPFF1[61]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(61));
    
    \RDATA_M_xhdl8[9]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9));
    
    \RDATA_M_int[44]\ : SLE
      port map(D => \RDATA_M_int_2[44]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[44]_net_1\);
    
    \WDATA_M_INPFF1[53]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(53), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[53]_net_1\);
    
    \RDATA_M_int[13]\ : SLE
      port map(D => \RDATA_M_int_2[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[13]_net_1\);
    
    \WDATA_M_INPFF1[14]\ : SLE
      port map(D => N_272_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[14]_net_1\);
    
    \WDATA_MI_xhdl22[36]\ : SLE
      port map(D => \WDATA_M_INPFF1[36]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(36));
    
    \RDATA_M_int[50]\ : SLE
      port map(D => \RDATA_M_int_2[50]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[50]_net_1\);
    
    \ARADDR_M_INPFF1[1]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(1));
    
    \WDATA_M_INPFF1[32]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(32), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[32]_net_1\);
    
    \RDATA_M_int[7]\ : SLE
      port map(D => \RDATA_M_int_2[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[7]_net_1\);
    
    \RDATA_M_int[5]\ : SLE
      port map(D => \RDATA_M_int_2[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[5]_net_1\);
    
    \L5.RDATA_M_xhdl8_3[62]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[62]_net_1\, Y
         => \RDATA_M_xhdl8_3[62]\);
    
    \WDATA_M_INPFF1[1]\ : SLE
      port map(D => N_136_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[1]_net_1\);
    
    \RDATA_M_int[60]\ : SLE
      port map(D => \RDATA_M_int_2[60]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[60]_net_1\);
    
    \RDATA_M_xhdl8[47]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[47]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47));
    
    \L5.RDATA_M_xhdl8_3[21]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[21]_net_1\, Y
         => \RDATA_M_xhdl8_3[21]\);
    
    \L5.RDATA_M_xhdl8_3[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[0]_net_1\, Y
         => \RDATA_M_xhdl8_3[0]\);
    
    \WDATA_MI_xhdl22[55]\ : SLE
      port map(D => \WDATA_M_INPFF1[55]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(55));
    
    \L5.RDATA_M_xhdl8_3[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[4]_net_1\, Y
         => \RDATA_M_xhdl8_3[4]\);
    
    \WDATA_MI_xhdl22[2]\ : SLE
      port map(D => \WDATA_M_INPFF1[2]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(2));
    
    \AWADDR_M_INPFF1[22]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(22));
    
    \WSTRB_MI_xhdl23[7]\ : SLE
      port map(D => \WSTRB_M_INPFF1[7]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(7));
    
    \WDATA_MI_xhdl22[49]\ : SLE
      port map(D => \WDATA_M_INPFF1[49]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(49));
    
    \AWADDR_M_INPFF1[17]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(17));
    
    \L5.RDATA_M_xhdl8_3[51]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[51]_net_1\, Y
         => \RDATA_M_xhdl8_3[51]\);
    
    \WSTRB_MI_xhdl23[2]\ : SLE
      port map(D => \WSTRB_M_INPFF1[2]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WSTRB_MI0(2));
    
    \WDATA_MI_xhdl22[8]\ : SLE
      port map(D => \WDATA_M_INPFF1[8]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(8));
    
    \L5.RDATA_M_xhdl8_3[47]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[47]_net_1\, Y
         => \RDATA_M_xhdl8_3[47]\);
    
    \L5.RDATA_M_xhdl8_3[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[12]_net_1\, Y
         => \RDATA_M_xhdl8_3[12]\);
    
    \AWLOCK_M_INPFF1[1]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, CLK => 
        SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWLOCK_MI0[1]\);
    
    \L5.RDATA_M_int_2[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(1), Y => 
        \RDATA_M_int_2[1]\);
    
    \WSTRB_M_INPFF1[0]\ : SLE
      port map(D => N_1445_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WSTRB_M_INPFF1[0]_net_1\);
    
    \WDATA_M_INPFF1[28]\ : SLE
      port map(D => N_197_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[28]_net_1\);
    
    \WDATA_M_INPFF1[19]\ : SLE
      port map(D => N_202_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[19]_net_1\);
    
    rdtrans_inprog : SLE
      port map(D => N_53, CLK => SDRCLK_c, EN => N_24, ALn => 
        MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rdtrans_inprog\);
    
    \L5.RDATA_M_xhdl8_3[28]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[28]_net_1\, Y
         => \RDATA_M_xhdl8_3[28]\);
    
    \RDATA_M_xhdl8[39]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[39]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39));
    
    \AWADDR_M_INPFF1[2]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(2));
    
    \RDATA_M_xhdl8[32]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[32]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32));
    
    \L5.RDATA_M_int_2[35]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(35), Y => 
        \RDATA_M_int_2[35]\);
    
    \WDATA_MI_xhdl22[40]\ : SLE
      port map(D => \WDATA_M_INPFF1[40]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(40));
    
    \L5.RDATA_M_xhdl8_3[58]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[58]_net_1\, Y
         => \RDATA_M_xhdl8_3[58]\);
    
    \L1.ARSIZE_M_INPFF1_2[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1), B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARREADY\, Y => 
        \ARSIZE_M_INPFF1_2[1]\);
    
    \L5.RDATA_M_int_2[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(16), Y => 
        \RDATA_M_int_2[16]\);
    
    \prev_ARADDR[26]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), CLK
         => SDRCLK_c, EN => N_28_i, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \prev_ARADDR[26]_net_1\);
    
    \WDATA_M_INPFF1[41]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(41), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[41]_net_1\);
    
    temp_xhdl44_2_i_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => N_34, B => \stall_trans\, Y => N_41);
    
    \RDATA_M_xhdl8[63]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[63]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63));
    
    \RDATA_M_xhdl8[36]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[36]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36));
    
    \RDATA_M_int[45]\ : SLE
      port map(D => \RDATA_M_int_2[45]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[45]_net_1\);
    
    \prev_ARADDR[27]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), CLK
         => SDRCLK_c, EN => N_28_i, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \prev_ARADDR[27]_net_1\);
    
    \L5.RDATA_M_int_2[55]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(55), Y => 
        \RDATA_M_int_2[55]\);
    
    \un1_rd_wdcntr_1_1.N_18_i\ : CFG4
      generic map(INIT => x"A965")

      port map(A => \rd_wdcntr[3]_net_1\, B => 
        \rd_wdcntr[2]_net_1\, C => N_37, D => N_36, Y => N_18_i);
    
    \L5.RDATA_M_int_2[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => RDATA_IM0(6), Y => 
        \RDATA_M_int_2[6]\);
    
    \L5.RDATA_M_xhdl8_3[46]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[46]_net_1\, Y
         => \RDATA_M_xhdl8_3[46]\);
    
    \WDATA_M_INPFF1[54]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_WDATA(54), CLK
         => SDRCLK_c, EN => \wready_m_xhdl2\, ALn => MSS_READY, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \WDATA_M_INPFF1[54]_net_1\);
    
    \WDATA_MI_xhdl22[15]\ : SLE
      port map(D => \WDATA_M_INPFF1[15]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(15));
    
    \RDATA_M_xhdl8[35]\ : SLE
      port map(D => \RDATA_M_xhdl8_3[35]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35));
    
    \ARADDR_M_INPFF1[18]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18), CLK
         => SDRCLK_c, EN => un2_arvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_MI0(18));
    
    \L5.RDATA_M_xhdl8_3[34]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \RREADY_MI0\, B => \RDATA_M_int[34]_net_1\, Y
         => \RDATA_M_xhdl8_3[34]\);
    
    \RDATA_M_int[41]\ : SLE
      port map(D => \RDATA_M_int_2[41]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[41]_net_1\);
    
    \WDATA_MI_xhdl22[35]\ : SLE
      port map(D => \WDATA_M_INPFF1[35]_net_1\, CLK => SDRCLK_c, 
        EN => \wready_m_xhdl2\, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => WDATA_MI0(35));
    
    \RDATA_M_int[53]\ : SLE
      port map(D => \RDATA_M_int_2[53]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_M_int[53]_net_1\);
    
    \WDATA_M_INPFF1[4]\ : SLE
      port map(D => N_133_i, CLK => SDRCLK_c, EN => 
        \wready_m_xhdl2\, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WDATA_M_INPFF1[4]_net_1\);
    
    \AWADDR_M_INPFF1[1]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1), CLK
         => SDRCLK_c, EN => un2_awvalid_m, ALn => MSS_READY, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_MI0(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_WA_ARBITER is

    port( AW_MASGNT_IC                         : out   std_logic_vector(3 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          AWLOCK_MI0_i_0                       : in    std_logic;
          m0_wr_end                            : in    std_logic;
          AW_REQ_MI0                           : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_WA_ARBITER;

architecture DEF_ARCH of axi_WA_ARBITER is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \wr_curr_state[12]_net_1\, \wr_curr_state_i[12]\, 
        \m0_lock_clear_write\, VCC_net_1, GND_net_1, N_128_i, 
        N_127_i, N_135_i, N_129_i, \wr_curr_state[8]_net_1\, 
        \wr_curr_state[7]_net_1\, \wr_curr_state[6]_net_1\, 
        N_110_i, \wr_curr_state[3]_net_1\, N_6, 
        \wr_curr_state[2]_net_1\, \wr_curr_state[1]_net_1\, 
        \wr_curr_state[0]_net_1\, \wr_curr_state[11]_net_1\, 
        \wr_curr_state_ns[1]_net_1\, \wr_curr_state[10]_net_1\, 
        \wr_curr_state_ns[2]\, \wr_curr_state[9]_net_1\, 
        \wr_curr_state_ns_0_a2_0[2]\, 
        \wr_curr_state_ns_o3[1]_net_1\, 
        \wr_curr_state_ns_i_i_a2_0[9]_net_1\, 
        \wr_curr_state_ns_0_o2[2]_net_1\ : std_logic;

begin 


    \AW_MASGNT_MI_xhdl1[1]\ : SLE
      port map(D => N_127_i, CLK => SDRCLK_c, EN => 
        \wr_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AW_MASGNT_IC(1));
    
    \wr_curr_state_ns_o3[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wr_curr_state[12]_net_1\, B => 
        \wr_curr_state[11]_net_1\, Y => 
        \wr_curr_state_ns_o3[1]_net_1\);
    
    \wr_curr_state[6]\ : SLE
      port map(D => N_110_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[6]_net_1\);
    
    m0_lock_clear_write : SLE
      port map(D => AWLOCK_MI0_i_0, CLK => SDRCLK_c, EN => 
        AW_REQ_MI0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \m0_lock_clear_write\);
    
    \wr_curr_state_RNO[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => m0_wr_end, B => \wr_curr_state[10]_net_1\, Y
         => N_110_i);
    
    \wr_curr_state_ns_0_o2[2]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => m0_wr_end, B => \m0_lock_clear_write\, C => 
        \wr_curr_state_ns_o3[1]_net_1\, D => 
        \wr_curr_state[3]_net_1\, Y => 
        \wr_curr_state_ns_0_o2[2]_net_1\);
    
    \wr_curr_state[0]\ : SLE
      port map(D => \wr_curr_state[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[0]_net_1\);
    
    \AW_MASGNT_MI_xhdl1_RNO[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wr_curr_state[3]_net_1\, B => 
        \wr_curr_state[10]_net_1\, Y => N_128_i);
    
    \wr_curr_state_ns_0_a2_0_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, B => 
        AW_REQ_MI0, Y => \wr_curr_state_ns_0_a2_0[2]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \wr_curr_state[10]\ : SLE
      port map(D => \wr_curr_state_ns[2]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[10]_net_1\);
    
    \wr_curr_state[9]\ : SLE
      port map(D => \wr_curr_state[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[9]_net_1\);
    
    \AW_MASGNT_MI_xhdl1_RNO[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wr_curr_state[0]_net_1\, B => 
        \wr_curr_state[7]_net_1\, Y => N_129_i);
    
    \AW_MASGNT_MI_xhdl1_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wr_curr_state[2]_net_1\, B => 
        \wr_curr_state[9]_net_1\, Y => N_127_i);
    
    \AW_MASGNT_MI_xhdl1[0]\ : SLE
      port map(D => N_128_i, CLK => SDRCLK_c, EN => 
        \wr_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AW_MASGNT_IC(0));
    
    \wr_curr_state_ns[1]\ : CFG3
      generic map(INIT => x"F4")

      port map(A => AW_REQ_MI0, B => 
        \wr_curr_state_ns_0_o2[2]_net_1\, C => 
        \wr_curr_state[6]_net_1\, Y => 
        \wr_curr_state_ns[1]_net_1\);
    
    \wr_curr_state_ns_0[2]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \wr_curr_state[10]_net_1\, B => m0_wr_end, C
         => \wr_curr_state_ns_0_a2_0[2]\, D => 
        \wr_curr_state_ns_0_o2[2]_net_1\, Y => 
        \wr_curr_state_ns[2]\);
    
    \wr_curr_state_ns_i_i_a2_0[9]\ : CFG4
      generic map(INIT => x"A800")

      port map(A => AW_REQ_MI0, B => \wr_curr_state[3]_net_1\, C
         => \wr_curr_state_ns_o3[1]_net_1\, D => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, Y => 
        \wr_curr_state_ns_i_i_a2_0[9]_net_1\);
    
    \wr_curr_state[2]\ : SLE
      port map(D => \wr_curr_state[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[2]_net_1\);
    
    \AW_MASGNT_MI_xhdl1_RNO[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \wr_curr_state[1]_net_1\, B => 
        \wr_curr_state[8]_net_1\, Y => N_135_i);
    
    \AW_MASGNT_MI_xhdl1[3]\ : SLE
      port map(D => N_129_i, CLK => SDRCLK_c, EN => 
        \wr_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AW_MASGNT_IC(3));
    
    \wr_curr_state_ns_i_i[9]\ : CFG4
      generic map(INIT => x"FF70")

      port map(A => \m0_lock_clear_write\, B => m0_wr_end, C => 
        \wr_curr_state[3]_net_1\, D => 
        \wr_curr_state_ns_i_i_a2_0[9]_net_1\, Y => N_6);
    
    \wr_curr_state[8]\ : SLE
      port map(D => \wr_curr_state[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[8]_net_1\);
    
    \AW_MASGNT_MI_xhdl1[2]\ : SLE
      port map(D => N_135_i, CLK => SDRCLK_c, EN => 
        \wr_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AW_MASGNT_IC(2));
    
    \wr_curr_state[1]\ : SLE
      port map(D => \wr_curr_state[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[1]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wr_curr_state_RNINP9[12]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wr_curr_state[12]_net_1\, Y => 
        \wr_curr_state_i[12]\);
    
    \wr_curr_state[12]\ : SLE
      port map(D => GND_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[12]_net_1\);
    
    \wr_curr_state[3]\ : SLE
      port map(D => N_6, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[3]_net_1\);
    
    \wr_curr_state[11]\ : SLE
      port map(D => \wr_curr_state_ns[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[11]_net_1\);
    
    \wr_curr_state[7]\ : SLE
      port map(D => \wr_curr_state[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wr_curr_state[7]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_wrmatrix_4Mto1S is

    port( AWSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1);
          AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWLOCK_MI0_i_0                       : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          MST_WRGNT_NUM_0                      : out   std_logic;
          m0_wr_end                            : in    std_logic;
          AWREADY_SI16                         : in    std_logic;
          AWVALID_MI0                          : in    std_logic;
          N_75_i                               : in    std_logic;
          AWVALID_IS16_gated                   : out   std_logic;
          AWREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_wrmatrix_4Mto1S;

architecture DEF_ARCH of axi_wrmatrix_4Mto1S is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component axi_WA_ARBITER
    port( AW_MASGNT_IC                         : out   std_logic_vector(3 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          AWLOCK_MI0_i_0                       : in    std_logic := 'U';
          m0_wr_end                            : in    std_logic := 'U';
          AW_REQ_MI0                           : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \AWSIZE_IS_int[0]_net_1\, VCC_net_1, 
        \AWSIZE_IS_int_2[0]\, GND_net_1, \AWSIZE_IS_int[1]_net_1\, 
        \AWSIZE_IS_int_2[1]\, \AWADDR_IS_int_xhdl7[17]_net_1\, 
        awaddr_is_int_xhdl74, \AWADDR_IS_int_xhdl7[18]_net_1\, 
        \AWADDR_IS_int_xhdl7[19]_net_1\, 
        \AWADDR_IS_int_xhdl7[20]_net_1\, 
        \AWADDR_IS_int_xhdl7[21]_net_1\, 
        \AWADDR_IS_int_xhdl7[22]_net_1\, 
        \AWADDR_IS_int_xhdl7[23]_net_1\, 
        \AWADDR_IS_int_xhdl7[26]_net_1\, 
        \AWADDR_IS_int_xhdl7[27]_net_1\, 
        \AWADDR_IS_int_xhdl7[2]_net_1\, 
        \AWADDR_IS_int_xhdl7[3]_net_1\, 
        \AWADDR_IS_int_xhdl7[4]_net_1\, 
        \AWADDR_IS_int_xhdl7[5]_net_1\, 
        \AWADDR_IS_int_xhdl7[6]_net_1\, 
        \AWADDR_IS_int_xhdl7[7]_net_1\, 
        \AWADDR_IS_int_xhdl7[8]_net_1\, 
        \AWADDR_IS_int_xhdl7[9]_net_1\, 
        \AWADDR_IS_int_xhdl7[10]_net_1\, 
        \AWADDR_IS_int_xhdl7[11]_net_1\, 
        \AWADDR_IS_int_xhdl7[12]_net_1\, 
        \AWADDR_IS_int_xhdl7[13]_net_1\, 
        \AWADDR_IS_int_xhdl7[14]_net_1\, 
        \AWADDR_IS_int_xhdl7[15]_net_1\, 
        \AWADDR_IS_int_xhdl7[16]_net_1\, 
        \AWADDR_IS_int_xhdl7[1]_net_1\, AWREADY_IM0_xhdl1_2, 
        \AWVALID_IS_int\, AWVALID_IS_int_2, \AW_REQ_MI0\, 
        \AW_MASGNT_IC[3]\, \AW_MASGNT_IC[2]\, \AW_MASGNT_IC[1]\, 
        \AW_MASGNT_IC[0]\ : std_logic;

    for all : axi_WA_ARBITER
	Use entity work.axi_WA_ARBITER(DEF_ARCH);
begin 


    \AWADDR_IS_int_xhdl7[22]\ : SLE
      port map(D => AWADDR_MI0(22), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[22]_net_1\);
    
    \AWADDR_IS_int_xhdl7[20]\ : SLE
      port map(D => AWADDR_MI0(20), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[20]_net_1\);
    
    \AWADDR_IS_xhdl6[14]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[14]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(14));
    
    \AWADDR_IS_int_xhdl7[27]\ : SLE
      port map(D => AWADDR_MI0(27), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[27]_net_1\);
    
    \L1.AWSIZE_IS_int_2[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => awaddr_is_int_xhdl74, B => AWSIZE_MI0(1), Y
         => \AWSIZE_IS_int_2[1]\);
    
    AW_REQ_MI0 : SLE
      port map(D => N_75_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \AW_REQ_MI0\);
    
    \AWADDR_IS_xhdl6[7]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[7]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(7));
    
    \AWADDR_IS_int_xhdl7[11]\ : SLE
      port map(D => AWADDR_MI0(11), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[11]_net_1\);
    
    \AWADDR_IS_int_xhdl7[9]\ : SLE
      port map(D => AWADDR_MI0(9), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[9]_net_1\);
    
    \AWADDR_IS_xhdl6[2]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[2]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(2));
    
    \AWADDR_IS_int_xhdl7[12]\ : SLE
      port map(D => AWADDR_MI0(12), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[12]_net_1\);
    
    \AWADDR_IS_int_xhdl7[10]\ : SLE
      port map(D => AWADDR_MI0(10), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[10]_net_1\);
    
    \AWSIZE_IS_int[0]\ : SLE
      port map(D => \AWSIZE_IS_int_2[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWSIZE_IS_int[0]_net_1\);
    
    \AWADDR_IS_int_xhdl7[17]\ : SLE
      port map(D => AWADDR_MI0(17), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[17]_net_1\);
    
    \AWADDR_IS_xhdl6[13]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[13]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(13));
    
    UWA_ARBITER : axi_WA_ARBITER
      port map(AW_MASGNT_IC(3) => \AW_MASGNT_IC[3]\, 
        AW_MASGNT_IC(2) => \AW_MASGNT_IC[2]\, AW_MASGNT_IC(1) => 
        \AW_MASGNT_IC[1]\, AW_MASGNT_IC(0) => \AW_MASGNT_IC[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, AWLOCK_MI0_i_0 => 
        AWLOCK_MI0_i_0, m0_wr_end => m0_wr_end, AW_REQ_MI0 => 
        \AW_REQ_MI0\, SDRCLK_c => SDRCLK_c, MSS_READY => 
        MSS_READY);
    
    AWVALID_IS_int : SLE
      port map(D => AWVALID_IS_int_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWVALID_IS_int\);
    
    AWVALID_IS_xhdl14 : SLE
      port map(D => \AWVALID_IS_int\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWVALID_IS16_gated);
    
    \AWADDR_IS_xhdl6[23]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[23]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(23));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \AWADDR_IS_xhdl6[11]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[11]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(11));
    
    \L1.AWVALID_IS_int_2\ : CFG2
      generic map(INIT => x"8")

      port map(A => awaddr_is_int_xhdl74, B => AWVALID_MI0, Y => 
        AWVALID_IS_int_2);
    
    \AWADDR_IS_xhdl6[12]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[12]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(12));
    
    \AWADDR_IS_xhdl6[10]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[10]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(10));
    
    \AWADDR_IS_xhdl6[21]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[21]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(21));
    
    \AWADDR_IS_xhdl6[17]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[17]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(17));
    
    \AWADDR_IS_int_xhdl7[7]\ : SLE
      port map(D => AWADDR_MI0(7), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[7]_net_1\);
    
    \AWADDR_IS_xhdl6[22]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[22]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(22));
    
    \AWADDR_IS_xhdl6[20]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[20]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(20));
    
    \AWADDR_IS_int_xhdl7[2]\ : SLE
      port map(D => AWADDR_MI0(2), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[2]_net_1\);
    
    \AWADDR_IS_xhdl6[27]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[27]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(27));
    
    \AWSIZE_IS_int[1]\ : SLE
      port map(D => \AWSIZE_IS_int_2[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWSIZE_IS_int[1]_net_1\);
    
    \AWADDR_IS_int_xhdl7[8]\ : SLE
      port map(D => AWADDR_MI0(8), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \AWADDR_IS_int_xhdl7[26]\ : SLE
      port map(D => AWADDR_MI0(26), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[26]_net_1\);
    
    \AWADDR_IS_xhdl6[6]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[6]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(6));
    
    \AWADDR_IS_xhdl6[4]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[4]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(4));
    
    \L1.awaddr_is_int_xhdl74\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \AW_MASGNT_IC[3]\, B => \AW_MASGNT_IC[2]\, C
         => \AW_MASGNT_IC[1]\, D => \AW_MASGNT_IC[0]\, Y => 
        awaddr_is_int_xhdl74);
    
    \AWADDR_IS_int_xhdl7[16]\ : SLE
      port map(D => AWADDR_MI0(16), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[16]_net_1\);
    
    AWREADY_IM0_xhdl1 : SLE
      port map(D => AWREADY_IM0_xhdl1_2, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWREADY_IM0);
    
    \AWADDR_IS_int_xhdl7[4]\ : SLE
      port map(D => AWADDR_MI0(4), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[4]_net_1\);
    
    \AWADDR_IS_int_xhdl7[1]\ : SLE
      port map(D => AWADDR_MI0(1), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[1]_net_1\);
    
    \AWADDR_IS_int_xhdl7[19]\ : SLE
      port map(D => AWADDR_MI0(19), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[19]_net_1\);
    
    \AWSIZE_IS_xhdl9[1]\ : SLE
      port map(D => \AWSIZE_IS_int[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWSIZE_IS16_gated(1));
    
    \L1.AWSIZE_IS_int_2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => awaddr_is_int_xhdl74, B => AWSIZE_MI0(0), Y
         => \AWSIZE_IS_int_2[0]\);
    
    \AWADDR_IS_int_xhdl7[18]\ : SLE
      port map(D => AWADDR_MI0(18), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[18]_net_1\);
    
    \AWADDR_IS_int_xhdl7[15]\ : SLE
      port map(D => AWADDR_MI0(15), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[15]_net_1\);
    
    \AWADDR_IS_xhdl6[5]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[5]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(5));
    
    \AWADDR_IS_int_xhdl7[3]\ : SLE
      port map(D => AWADDR_MI0(3), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[3]_net_1\);
    
    \MST_WRGNT_NUM_xhdl16[0]\ : SLE
      port map(D => awaddr_is_int_xhdl74, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        MST_WRGNT_NUM_0);
    
    \AWADDR_IS_xhdl6[9]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[9]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(9));
    
    \AWADDR_IS_xhdl6[8]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[8]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(8));
    
    \L1.AWREADY_IM0_xhdl1_2\ : CFG2
      generic map(INIT => x"4")

      port map(A => AWREADY_SI16, B => awaddr_is_int_xhdl74, Y
         => AWREADY_IM0_xhdl1_2);
    
    \AWSIZE_IS_xhdl9[0]\ : SLE
      port map(D => \AWSIZE_IS_int[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        AWSIZE_IS16_gated(0));
    
    \AWADDR_IS_xhdl6[16]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[16]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(16));
    
    \AWADDR_IS_int_xhdl7[14]\ : SLE
      port map(D => AWADDR_MI0(14), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[14]_net_1\);
    
    \AWADDR_IS_int_xhdl7[23]\ : SLE
      port map(D => AWADDR_MI0(23), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[23]_net_1\);
    
    \AWADDR_IS_xhdl6[1]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[1]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(1));
    
    \AWADDR_IS_xhdl6[19]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[19]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(19));
    
    \AWADDR_IS_xhdl6[26]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[26]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(26));
    
    \AWADDR_IS_xhdl6[18]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[18]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(18));
    
    \AWADDR_IS_int_xhdl7[6]\ : SLE
      port map(D => AWADDR_MI0(6), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[6]_net_1\);
    
    \AWADDR_IS_xhdl6[15]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[15]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(15));
    
    \AWADDR_IS_int_xhdl7[13]\ : SLE
      port map(D => AWADDR_MI0(13), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[13]_net_1\);
    
    \AWADDR_IS_xhdl6[3]\ : SLE
      port map(D => \AWADDR_IS_int_xhdl7[3]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => AWADDR_IS16_gated(3));
    
    \AWADDR_IS_int_xhdl7[5]\ : SLE
      port map(D => AWADDR_MI0(5), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[5]_net_1\);
    
    \AWADDR_IS_int_xhdl7[21]\ : SLE
      port map(D => AWADDR_MI0(21), CLK => SDRCLK_c, EN => 
        awaddr_is_int_xhdl74, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \AWADDR_IS_int_xhdl7[21]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_wa_channel is

    port( AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1);
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          MST_WRGNT_NUM_0                      : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          AWLOCK_MI0_i_0                       : in    std_logic;
          MSS_READY                            : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          AWREADY_IM0                          : out   std_logic;
          AWVALID_IS16_gated                   : out   std_logic;
          N_75_i                               : in    std_logic;
          AWVALID_MI0                          : in    std_logic;
          AWREADY_SI16                         : in    std_logic;
          m0_wr_end                            : in    std_logic
        );

end axi_wa_channel;

architecture DEF_ARCH of axi_wa_channel is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component axi_wrmatrix_4Mto1S
    port( AWSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWLOCK_MI0_i_0                       : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          MST_WRGNT_NUM_0                      : out   std_logic;
          m0_wr_end                            : in    std_logic := 'U';
          AWREADY_SI16                         : in    std_logic := 'U';
          AWVALID_MI0                          : in    std_logic := 'U';
          N_75_i                               : in    std_logic := 'U';
          AWVALID_IS16_gated                   : out   std_logic;
          AWREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : axi_wrmatrix_4Mto1S
	Use entity work.axi_wrmatrix_4Mto1S(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \L1.inst_wrmatrix_4Mto1S\ : axi_wrmatrix_4Mto1S
      port map(AWSIZE_MI0(1) => AWSIZE_MI0(1), AWSIZE_MI0(0) => 
        AWSIZE_MI0(0), AWADDR_IS16_gated(27) => 
        AWADDR_IS16_gated(27), AWADDR_IS16_gated(26) => 
        AWADDR_IS16_gated(26), AWADDR_IS16_gated(25) => nc2, 
        AWADDR_IS16_gated(24) => nc4, AWADDR_IS16_gated(23) => 
        AWADDR_IS16_gated(23), AWADDR_IS16_gated(22) => 
        AWADDR_IS16_gated(22), AWADDR_IS16_gated(21) => 
        AWADDR_IS16_gated(21), AWADDR_IS16_gated(20) => 
        AWADDR_IS16_gated(20), AWADDR_IS16_gated(19) => 
        AWADDR_IS16_gated(19), AWADDR_IS16_gated(18) => 
        AWADDR_IS16_gated(18), AWADDR_IS16_gated(17) => 
        AWADDR_IS16_gated(17), AWADDR_IS16_gated(16) => 
        AWADDR_IS16_gated(16), AWADDR_IS16_gated(15) => 
        AWADDR_IS16_gated(15), AWADDR_IS16_gated(14) => 
        AWADDR_IS16_gated(14), AWADDR_IS16_gated(13) => 
        AWADDR_IS16_gated(13), AWADDR_IS16_gated(12) => 
        AWADDR_IS16_gated(12), AWADDR_IS16_gated(11) => 
        AWADDR_IS16_gated(11), AWADDR_IS16_gated(10) => 
        AWADDR_IS16_gated(10), AWADDR_IS16_gated(9) => 
        AWADDR_IS16_gated(9), AWADDR_IS16_gated(8) => 
        AWADDR_IS16_gated(8), AWADDR_IS16_gated(7) => 
        AWADDR_IS16_gated(7), AWADDR_IS16_gated(6) => 
        AWADDR_IS16_gated(6), AWADDR_IS16_gated(5) => 
        AWADDR_IS16_gated(5), AWADDR_IS16_gated(4) => 
        AWADDR_IS16_gated(4), AWADDR_IS16_gated(3) => 
        AWADDR_IS16_gated(3), AWADDR_IS16_gated(2) => 
        AWADDR_IS16_gated(2), AWADDR_IS16_gated(1) => 
        AWADDR_IS16_gated(1), AWADDR_MI0(27) => AWADDR_MI0(27), 
        AWADDR_MI0(26) => AWADDR_MI0(26), AWADDR_MI0(25) => nc3, 
        AWADDR_MI0(24) => nc1, AWADDR_MI0(23) => AWADDR_MI0(23), 
        AWADDR_MI0(22) => AWADDR_MI0(22), AWADDR_MI0(21) => 
        AWADDR_MI0(21), AWADDR_MI0(20) => AWADDR_MI0(20), 
        AWADDR_MI0(19) => AWADDR_MI0(19), AWADDR_MI0(18) => 
        AWADDR_MI0(18), AWADDR_MI0(17) => AWADDR_MI0(17), 
        AWADDR_MI0(16) => AWADDR_MI0(16), AWADDR_MI0(15) => 
        AWADDR_MI0(15), AWADDR_MI0(14) => AWADDR_MI0(14), 
        AWADDR_MI0(13) => AWADDR_MI0(13), AWADDR_MI0(12) => 
        AWADDR_MI0(12), AWADDR_MI0(11) => AWADDR_MI0(11), 
        AWADDR_MI0(10) => AWADDR_MI0(10), AWADDR_MI0(9) => 
        AWADDR_MI0(9), AWADDR_MI0(8) => AWADDR_MI0(8), 
        AWADDR_MI0(7) => AWADDR_MI0(7), AWADDR_MI0(6) => 
        AWADDR_MI0(6), AWADDR_MI0(5) => AWADDR_MI0(5), 
        AWADDR_MI0(4) => AWADDR_MI0(4), AWADDR_MI0(3) => 
        AWADDR_MI0(3), AWADDR_MI0(2) => AWADDR_MI0(2), 
        AWADDR_MI0(1) => AWADDR_MI0(1), AWSIZE_IS16_gated(1) => 
        AWSIZE_IS16_gated(1), AWSIZE_IS16_gated(0) => 
        AWSIZE_IS16_gated(0), AWLOCK_MI0_i_0 => AWLOCK_MI0_i_0, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, MST_WRGNT_NUM_0 => 
        MST_WRGNT_NUM_0, m0_wr_end => m0_wr_end, AWREADY_SI16 => 
        AWREADY_SI16, AWVALID_MI0 => AWVALID_MI0, N_75_i => 
        N_75_i, AWVALID_IS16_gated => AWVALID_IS16_gated, 
        AWREADY_IM0 => AWREADY_IM0, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_wd_channel is

    port( WDATA_MI0         : in    std_logic_vector(63 downto 0);
          WSTRB_MI0         : in    std_logic_vector(7 downto 0);
          WDATA_IS16_gated  : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated  : out   std_logic_vector(7 downto 0);
          MST_WRGNT_NUM_0   : in    std_logic;
          WREADY_SI16       : in    std_logic;
          WVALID_MI0        : in    std_logic;
          WVALID_IS16_gated : out   std_logic;
          WREADY_IM0        : out   std_logic;
          SDRCLK_c          : in    std_logic;
          MSS_READY         : in    std_logic
        );

end axi_wd_channel;

architecture DEF_ARCH of axi_wd_channel is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \MST_GNT_NUM_r[0]_net_1\, VCC_net_1, GND_net_1, 
        \WDATA_IS_xhdl6_3[51]_net_1\, 
        \WDATA_IS_xhdl6_3[52]_net_1\, 
        \WDATA_IS_xhdl6_3[53]_net_1\, 
        \WDATA_IS_xhdl6_3[54]_net_1\, 
        \WDATA_IS_xhdl6_3[55]_net_1\, 
        \WDATA_IS_xhdl6_3[56]_net_1\, 
        \WDATA_IS_xhdl6_3[57]_net_1\, 
        \WDATA_IS_xhdl6_3[58]_net_1\, 
        \WDATA_IS_xhdl6_3[59]_net_1\, 
        \WDATA_IS_xhdl6_3[60]_net_1\, 
        \WDATA_IS_xhdl6_3[61]_net_1\, 
        \WDATA_IS_xhdl6_3[62]_net_1\, 
        \WDATA_IS_xhdl6_3[63]_net_1\, 
        \WDATA_IS_xhdl6_3[36]_net_1\, 
        \WDATA_IS_xhdl6_3[37]_net_1\, 
        \WDATA_IS_xhdl6_3[38]_net_1\, 
        \WDATA_IS_xhdl6_3[39]_net_1\, 
        \WDATA_IS_xhdl6_3[40]_net_1\, 
        \WDATA_IS_xhdl6_3[41]_net_1\, 
        \WDATA_IS_xhdl6_3[42]_net_1\, 
        \WDATA_IS_xhdl6_3[43]_net_1\, 
        \WDATA_IS_xhdl6_3[44]_net_1\, 
        \WDATA_IS_xhdl6_3[45]_net_1\, 
        \WDATA_IS_xhdl6_3[46]_net_1\, 
        \WDATA_IS_xhdl6_3[47]_net_1\, 
        \WDATA_IS_xhdl6_3[48]_net_1\, 
        \WDATA_IS_xhdl6_3[49]_net_1\, 
        \WDATA_IS_xhdl6_3[50]_net_1\, 
        \WDATA_IS_xhdl6_3[21]_net_1\, 
        \WDATA_IS_xhdl6_3[22]_net_1\, 
        \WDATA_IS_xhdl6_3[23]_net_1\, 
        \WDATA_IS_xhdl6_3[24]_net_1\, 
        \WDATA_IS_xhdl6_3[25]_net_1\, 
        \WDATA_IS_xhdl6_3[26]_net_1\, 
        \WDATA_IS_xhdl6_3[27]_net_1\, 
        \WDATA_IS_xhdl6_3[28]_net_1\, 
        \WDATA_IS_xhdl6_3[29]_net_1\, 
        \WDATA_IS_xhdl6_3[30]_net_1\, 
        \WDATA_IS_xhdl6_3[31]_net_1\, 
        \WDATA_IS_xhdl6_3[32]_net_1\, 
        \WDATA_IS_xhdl6_3[33]_net_1\, 
        \WDATA_IS_xhdl6_3[34]_net_1\, 
        \WDATA_IS_xhdl6_3[35]_net_1\, \WDATA_IS_xhdl6_3[6]_net_1\, 
        \WDATA_IS_xhdl6_3[7]_net_1\, \WDATA_IS_xhdl6_3[8]_net_1\, 
        \WDATA_IS_xhdl6_3[9]_net_1\, \WDATA_IS_xhdl6_3[10]_net_1\, 
        \WDATA_IS_xhdl6_3[11]_net_1\, 
        \WDATA_IS_xhdl6_3[12]_net_1\, 
        \WDATA_IS_xhdl6_3[13]_net_1\, 
        \WDATA_IS_xhdl6_3[14]_net_1\, 
        \WDATA_IS_xhdl6_3[15]_net_1\, 
        \WDATA_IS_xhdl6_3[16]_net_1\, 
        \WDATA_IS_xhdl6_3[17]_net_1\, 
        \WDATA_IS_xhdl6_3[18]_net_1\, 
        \WDATA_IS_xhdl6_3[19]_net_1\, 
        \WDATA_IS_xhdl6_3[20]_net_1\, \WSTRB_IS_xhdl7_3[0]_net_1\, 
        \WSTRB_IS_xhdl7_3[1]_net_1\, \WSTRB_IS_xhdl7_3[2]_net_1\, 
        \WSTRB_IS_xhdl7_3[3]_net_1\, \WSTRB_IS_xhdl7_3[4]_net_1\, 
        \WSTRB_IS_xhdl7_3[5]_net_1\, \WSTRB_IS_xhdl7_3[6]_net_1\, 
        \WSTRB_IS_xhdl7_3[7]_net_1\, \WDATA_IS_xhdl6_3[0]_net_1\, 
        \WDATA_IS_xhdl6_3[1]_net_1\, \WDATA_IS_xhdl6_3[2]_net_1\, 
        \WDATA_IS_xhdl6_3[3]_net_1\, \WDATA_IS_xhdl6_3[4]_net_1\, 
        \WDATA_IS_xhdl6_3[5]_net_1\, wready_im0_int_xhdl15_1, 
        \WVALID_IS_xhdl9_2\ : std_logic;

begin 


    \WDATA_IS_xhdl6[50]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[50]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(50));
    
    \WDATA_IS_xhdl6_3[39]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(39), Y => 
        \WDATA_IS_xhdl6_3[39]_net_1\);
    
    \WSTRB_IS_xhdl7[6]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[6]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(6));
    
    \WDATA_IS_xhdl6_3[23]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(23), Y => 
        \WDATA_IS_xhdl6_3[23]_net_1\);
    
    \WDATA_IS_xhdl6_3[14]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(14), Y => 
        \WDATA_IS_xhdl6_3[14]_net_1\);
    
    \WDATA_IS_xhdl6[62]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[62]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(62));
    
    \WDATA_IS_xhdl6[0]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[0]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(0));
    
    \WDATA_IS_xhdl6[48]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[48]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(48));
    
    \WSTRB_IS_xhdl7_3[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(5), Y => 
        \WSTRB_IS_xhdl7_3[5]_net_1\);
    
    \WDATA_IS_xhdl6_3[16]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(16), Y => 
        \WDATA_IS_xhdl6_3[16]_net_1\);
    
    \WDATA_IS_xhdl6_3[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(15), Y => 
        \WDATA_IS_xhdl6_3[15]_net_1\);
    
    \WDATA_IS_xhdl6_3[60]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(60), Y => 
        \WDATA_IS_xhdl6_3[60]_net_1\);
    
    \WDATA_IS_xhdl6[42]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[42]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(42));
    
    \WDATA_IS_xhdl6[58]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[58]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(58));
    
    \WDATA_IS_xhdl6[17]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[17]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(17));
    
    \WSTRB_IS_xhdl7_3[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(3), Y => 
        \WSTRB_IS_xhdl7_3[3]_net_1\);
    
    \WDATA_IS_xhdl6[52]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[52]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(52));
    
    \WDATA_IS_xhdl6[19]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[19]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(19));
    
    \WDATA_IS_xhdl6_3[48]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(48), Y => 
        \WDATA_IS_xhdl6_3[48]_net_1\);
    
    \WDATA_IS_xhdl6[37]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[37]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(37));
    
    \WSTRB_IS_xhdl7[3]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[3]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(3));
    
    \WDATA_IS_xhdl6[39]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[39]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(39));
    
    \WDATA_IS_xhdl6_3[28]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(28), Y => 
        \WDATA_IS_xhdl6_3[28]_net_1\);
    
    \WDATA_IS_xhdl6_3[37]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(37), Y => 
        \WDATA_IS_xhdl6_3[37]_net_1\);
    
    \WDATA_IS_xhdl6[14]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[14]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(14));
    
    \WDATA_IS_xhdl6_3[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(9), Y => 
        \WDATA_IS_xhdl6_3[9]_net_1\);
    
    \WDATA_IS_xhdl6_3[44]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(44), Y => 
        \WDATA_IS_xhdl6_3[44]_net_1\);
    
    \WDATA_IS_xhdl6[11]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[11]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(11));
    
    WVALID_IS_xhdl9_2 : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WVALID_MI0, Y => 
        \WVALID_IS_xhdl9_2\);
    
    \WDATA_IS_xhdl6[34]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[34]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(34));
    
    \WDATA_IS_xhdl6_3[46]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(46), Y => 
        \WDATA_IS_xhdl6_3[46]_net_1\);
    
    \WDATA_IS_xhdl6_3[45]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(45), Y => 
        \WDATA_IS_xhdl6_3[45]_net_1\);
    
    \WDATA_IS_xhdl6_3[24]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(24), Y => 
        \WDATA_IS_xhdl6_3[24]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \WDATA_IS_xhdl6[31]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[31]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(31));
    
    \WDATA_IS_xhdl6[8]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[8]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(8));
    
    \WDATA_IS_xhdl6_3[26]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(26), Y => 
        \WDATA_IS_xhdl6_3[26]_net_1\);
    
    \WDATA_IS_xhdl6_3[25]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(25), Y => 
        \WDATA_IS_xhdl6_3[25]_net_1\);
    
    \WDATA_IS_xhdl6_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(0), Y => 
        \WDATA_IS_xhdl6_3[0]_net_1\);
    
    \WDATA_IS_xhdl6_3[50]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(50), Y => 
        \WDATA_IS_xhdl6_3[50]_net_1\);
    
    \WDATA_IS_xhdl6_3[32]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(32), Y => 
        \WDATA_IS_xhdl6_3[32]_net_1\);
    
    \WDATA_IS_xhdl6[23]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[23]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(23));
    
    \WDATA_IS_xhdl6_3[31]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(31), Y => 
        \WDATA_IS_xhdl6_3[31]_net_1\);
    
    \WDATA_IS_xhdl6_3[59]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(59), Y => 
        \WDATA_IS_xhdl6_3[59]_net_1\);
    
    \WDATA_IS_xhdl6[10]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[10]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(10));
    
    \WDATA_IS_xhdl6_3[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(2), Y => 
        \WDATA_IS_xhdl6_3[2]_net_1\);
    
    \WDATA_IS_xhdl6[1]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(1));
    
    \WDATA_IS_xhdl6_3[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(1), Y => 
        \WDATA_IS_xhdl6_3[1]_net_1\);
    
    \WSTRB_IS_xhdl7_3[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(7), Y => 
        \WSTRB_IS_xhdl7_3[7]_net_1\);
    
    \WDATA_IS_xhdl6_3[62]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(62), Y => 
        \WDATA_IS_xhdl6_3[62]_net_1\);
    
    \WDATA_IS_xhdl6[30]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[30]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(30));
    
    \WDATA_IS_xhdl6[63]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[63]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(63));
    
    \WDATA_IS_xhdl6_3[61]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(61), Y => 
        \WDATA_IS_xhdl6_3[61]_net_1\);
    
    \WDATA_IS_xhdl6[18]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[18]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(18));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \WDATA_IS_xhdl6_3[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(10), Y => 
        \WDATA_IS_xhdl6_3[10]_net_1\);
    
    \WDATA_IS_xhdl6[43]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[43]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(43));
    
    \WDATA_IS_xhdl6[12]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[12]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(12));
    
    \WSTRB_IS_xhdl7_3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(6), Y => 
        \WSTRB_IS_xhdl7_3[6]_net_1\);
    
    \WDATA_IS_xhdl6[38]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[38]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(38));
    
    \WDATA_IS_xhdl6[53]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[53]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(53));
    
    \WDATA_IS_xhdl6[32]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[32]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(32));
    
    \WDATA_IS_xhdl6[6]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[6]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(6));
    
    \WSTRB_IS_xhdl7_3[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(1), Y => 
        \WSTRB_IS_xhdl7_3[1]_net_1\);
    
    \WDATA_IS_xhdl6_3[19]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(19), Y => 
        \WDATA_IS_xhdl6_3[19]_net_1\);
    
    \WDATA_IS_xhdl6_3[57]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(57), Y => 
        \WDATA_IS_xhdl6_3[57]_net_1\);
    
    \WDATA_IS_xhdl6_3[33]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(33), Y => 
        \WDATA_IS_xhdl6_3[33]_net_1\);
    
    WVALID_IS_xhdl9 : SLE
      port map(D => \WVALID_IS_xhdl9_2\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WVALID_IS16_gated);
    
    \WSTRB_IS_xhdl7_3[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(2), Y => 
        \WSTRB_IS_xhdl7_3[2]_net_1\);
    
    \WDATA_IS_xhdl6[9]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[9]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(9));
    
    \WDATA_IS_xhdl6[25]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[25]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(25));
    
    \WDATA_IS_xhdl6_3[63]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(63), Y => 
        \WDATA_IS_xhdl6_3[63]_net_1\);
    
    \WDATA_IS_xhdl6_3[38]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(38), Y => 
        \WDATA_IS_xhdl6_3[38]_net_1\);
    
    \WDATA_IS_xhdl6_3[40]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(40), Y => 
        \WDATA_IS_xhdl6_3[40]_net_1\);
    
    \WDATA_IS_xhdl6_3[17]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(17), Y => 
        \WDATA_IS_xhdl6_3[17]_net_1\);
    
    \WDATA_IS_xhdl6[7]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[7]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(7));
    
    \WDATA_IS_xhdl6[26]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[26]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(26));
    
    \WDATA_IS_xhdl6_3[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(20), Y => 
        \WDATA_IS_xhdl6_3[20]_net_1\);
    
    \WDATA_IS_xhdl6_3[52]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(52), Y => 
        \WDATA_IS_xhdl6_3[52]_net_1\);
    
    \WDATA_IS_xhdl6[3]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[3]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(3));
    
    \WSTRB_IS_xhdl7[0]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[0]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(0));
    
    \WDATA_IS_xhdl6_3[51]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(51), Y => 
        \WDATA_IS_xhdl6_3[51]_net_1\);
    
    \WDATA_IS_xhdl6_3[49]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(49), Y => 
        \WDATA_IS_xhdl6_3[49]_net_1\);
    
    \WDATA_IS_xhdl6[45]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[45]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(45));
    
    \WDATA_IS_xhdl6_3[29]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(29), Y => 
        \WDATA_IS_xhdl6_3[29]_net_1\);
    
    \WDATA_IS_xhdl6_3[34]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(34), Y => 
        \WDATA_IS_xhdl6_3[34]_net_1\);
    
    \WDATA_IS_xhdl6[55]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[55]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(55));
    
    \WDATA_IS_xhdl6[27]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[27]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(27));
    
    \WDATA_IS_xhdl6_3[36]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(36), Y => 
        \WDATA_IS_xhdl6_3[36]_net_1\);
    
    \WDATA_IS_xhdl6_3[35]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(35), Y => 
        \WDATA_IS_xhdl6_3[35]_net_1\);
    
    \L1.wready_im0_int_xhdl15_1\ : CFG2
      generic map(INIT => x"8")

      port map(A => WREADY_SI16, B => \MST_GNT_NUM_r[0]_net_1\, Y
         => wready_im0_int_xhdl15_1);
    
    \WDATA_IS_xhdl6[29]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[29]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(29));
    
    \WDATA_IS_xhdl6[46]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[46]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(46));
    
    \WSTRB_IS_xhdl7_3[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(4), Y => 
        \WSTRB_IS_xhdl7_3[4]_net_1\);
    
    \WDATA_IS_xhdl6_3[12]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(12), Y => 
        \WDATA_IS_xhdl6_3[12]_net_1\);
    
    \WDATA_IS_xhdl6[56]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[56]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(56));
    
    \WDATA_IS_xhdl6_3[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(7), Y => 
        \WDATA_IS_xhdl6_3[7]_net_1\);
    
    \WDATA_IS_xhdl6_3[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(11), Y => 
        \WDATA_IS_xhdl6_3[11]_net_1\);
    
    \WDATA_IS_xhdl6_3[47]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(47), Y => 
        \WDATA_IS_xhdl6_3[47]_net_1\);
    
    \WSTRB_IS_xhdl7[5]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[5]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(5));
    
    \WDATA_IS_xhdl6[13]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[13]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(13));
    
    \WDATA_IS_xhdl6_3[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(4), Y => 
        \WDATA_IS_xhdl6_3[4]_net_1\);
    
    \WDATA_IS_xhdl6_3[27]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(27), Y => 
        \WDATA_IS_xhdl6_3[27]_net_1\);
    
    \WDATA_IS_xhdl6_3[53]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(53), Y => 
        \WDATA_IS_xhdl6_3[53]_net_1\);
    
    \WDATA_IS_xhdl6[47]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[47]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(47));
    
    \WDATA_IS_xhdl6[33]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[33]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(33));
    
    \WDATA_IS_xhdl6[4]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[4]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(4));
    
    \WDATA_IS_xhdl6[24]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[24]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(24));
    
    \WDATA_IS_xhdl6[49]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[49]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(49));
    
    \WDATA_IS_xhdl6[57]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[57]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(57));
    
    \WDATA_IS_xhdl6[21]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[21]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(21));
    
    \WDATA_IS_xhdl6[5]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[5]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(5));
    
    \WDATA_IS_xhdl6[59]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[59]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(59));
    
    WREADY_IM0_xhdl1 : SLE
      port map(D => wready_im0_int_xhdl15_1, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WREADY_IM0);
    
    \WSTRB_IS_xhdl7[2]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[2]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(2));
    
    \WDATA_IS_xhdl6_3[58]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(58), Y => 
        \WDATA_IS_xhdl6_3[58]_net_1\);
    
    \WSTRB_IS_xhdl7[7]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[7]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(7));
    
    \WDATA_IS_xhdl6_3[42]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(42), Y => 
        \WDATA_IS_xhdl6_3[42]_net_1\);
    
    \WDATA_IS_xhdl6_3[13]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(13), Y => 
        \WDATA_IS_xhdl6_3[13]_net_1\);
    
    \WDATA_IS_xhdl6[44]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[44]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(44));
    
    \WDATA_IS_xhdl6[61]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[61]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(61));
    
    \WDATA_IS_xhdl6_3[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(5), Y => 
        \WDATA_IS_xhdl6_3[5]_net_1\);
    
    \WDATA_IS_xhdl6_3[41]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(41), Y => 
        \WDATA_IS_xhdl6_3[41]_net_1\);
    
    \WDATA_IS_xhdl6[54]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[54]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(54));
    
    \WDATA_IS_xhdl6[41]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[41]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(41));
    
    \WDATA_IS_xhdl6_3[22]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(22), Y => 
        \WDATA_IS_xhdl6_3[22]_net_1\);
    
    \MST_GNT_NUM_r[0]\ : SLE
      port map(D => MST_WRGNT_NUM_0, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MST_GNT_NUM_r[0]_net_1\);
    
    \WDATA_IS_xhdl6_3[21]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(21), Y => 
        \WDATA_IS_xhdl6_3[21]_net_1\);
    
    \WDATA_IS_xhdl6[51]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[51]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(51));
    
    \WDATA_IS_xhdl6[20]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[20]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(20));
    
    \WDATA_IS_xhdl6_3[54]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(54), Y => 
        \WDATA_IS_xhdl6_3[54]_net_1\);
    
    \WDATA_IS_xhdl6_3[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(8), Y => 
        \WDATA_IS_xhdl6_3[8]_net_1\);
    
    \WDATA_IS_xhdl6[2]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[2]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(2));
    
    \WDATA_IS_xhdl6_3[18]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(18), Y => 
        \WDATA_IS_xhdl6_3[18]_net_1\);
    
    \WDATA_IS_xhdl6_3[56]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(56), Y => 
        \WDATA_IS_xhdl6_3[56]_net_1\);
    
    \WDATA_IS_xhdl6[15]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[15]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(15));
    
    \WDATA_IS_xhdl6_3[55]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(55), Y => 
        \WDATA_IS_xhdl6_3[55]_net_1\);
    
    \WDATA_IS_xhdl6[28]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[28]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(28));
    
    \WDATA_IS_xhdl6[35]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[35]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(35));
    
    \WDATA_IS_xhdl6[22]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[22]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(22));
    
    \WDATA_IS_xhdl6_3[30]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(30), Y => 
        \WDATA_IS_xhdl6_3[30]_net_1\);
    
    \WDATA_IS_xhdl6[60]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[60]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(60));
    
    \WSTRB_IS_xhdl7[4]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[4]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(4));
    
    \WDATA_IS_xhdl6_3[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(3), Y => 
        \WDATA_IS_xhdl6_3[3]_net_1\);
    
    \WDATA_IS_xhdl6[16]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[16]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(16));
    
    \WSTRB_IS_xhdl7[1]\ : SLE
      port map(D => \WSTRB_IS_xhdl7_3[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WSTRB_IS16_gated(1));
    
    \WDATA_IS_xhdl6[40]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[40]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(40));
    
    \WDATA_IS_xhdl6_3[43]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(43), Y => 
        \WDATA_IS_xhdl6_3[43]_net_1\);
    
    \WSTRB_IS_xhdl7_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WSTRB_MI0(0), Y => 
        \WSTRB_IS_xhdl7_3[0]_net_1\);
    
    \WDATA_IS_xhdl6_3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => MST_WRGNT_NUM_0, B => WDATA_MI0(6), Y => 
        \WDATA_IS_xhdl6_3[6]_net_1\);
    
    \WDATA_IS_xhdl6[36]\ : SLE
      port map(D => \WDATA_IS_xhdl6_3[36]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        WDATA_IS16_gated(36));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_RA_ARBITER is

    port( AR_MASGNT_IC                         : out   std_logic_vector(3 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          ARLOCK_MI0_i_0                       : in    std_logic;
          m0_rd_end                            : in    std_logic;
          AR_REQ_MI0                           : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_RA_ARBITER;

architecture DEF_ARCH of axi_RA_ARBITER is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \rd_curr_state[12]_net_1\, \rd_curr_state_i[12]\, 
        \m0_lock_clear_read\, VCC_net_1, GND_net_1, N_142_i, 
        N_165_i, N_163_i, N_164_i, \rd_curr_state[9]_net_1\, 
        \rd_curr_state[8]_net_1\, \rd_curr_state[7]_net_1\, 
        \rd_curr_state_ns[6]\, \rd_curr_state[3]_net_1\, N_134_i, 
        \rd_curr_state[2]_net_1\, \rd_curr_state[1]_net_1\, 
        \rd_curr_state[0]_net_1\, \rd_curr_state[13]_net_1\, 
        \rd_curr_state_ns[0]\, \rd_curr_state_ns[1]_net_1\, 
        \rd_curr_state[11]_net_1\, \rd_curr_state_ns[2]_net_1\, 
        \rd_curr_state[10]_net_1\, N_150, N_152, N_158, N_151, 
        N_149, \rd_curr_state_ns_i_0[10]_net_1\ : std_logic;

begin 


    \AR_MASGNT_MI_xhdl1_RNO[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \rd_curr_state[0]_net_1\, B => 
        \rd_curr_state[8]_net_1\, Y => N_164_i);
    
    \rd_curr_state_RNINC3B[12]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rd_curr_state[12]_net_1\, Y => 
        \rd_curr_state_i[12]\);
    
    \rd_curr_state_ns_o2[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \rd_curr_state[11]_net_1\, B => N_150, C => 
        \rd_curr_state[12]_net_1\, Y => N_152);
    
    \rd_curr_state_ns_a2[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => AR_REQ_MI0, B => \rd_curr_state[12]_net_1\, Y
         => \rd_curr_state_ns[0]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \rd_curr_state[11]\ : SLE
      port map(D => \rd_curr_state_ns[2]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[11]_net_1\);
    
    \rd_curr_state[2]\ : SLE
      port map(D => \rd_curr_state[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[2]_net_1\);
    
    \rd_curr_state[12]\ : SLE
      port map(D => \rd_curr_state_ns[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[12]_net_1\);
    
    \rd_curr_state_ns_o2[1]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => \m0_lock_clear_read\, B => 
        \rd_curr_state[13]_net_1\, C => m0_rd_end, D => 
        \rd_curr_state[3]_net_1\, Y => N_150);
    
    \AR_MASGNT_MI_xhdl1_RNO[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \rd_curr_state[2]_net_1\, B => 
        \rd_curr_state[10]_net_1\, Y => N_165_i);
    
    \rd_curr_state_ns[1]\ : CFG3
      generic map(INIT => x"CE")

      port map(A => N_150, B => \rd_curr_state[7]_net_1\, C => 
        AR_REQ_MI0, Y => \rd_curr_state_ns[1]_net_1\);
    
    \rd_curr_state[7]\ : SLE
      port map(D => \rd_curr_state_ns[6]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[7]_net_1\);
    
    \rd_curr_state[3]\ : SLE
      port map(D => N_134_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[3]_net_1\);
    
    \rd_curr_state_ns_i_o3[10]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \rd_curr_state[11]_net_1\, B => 
        \rd_curr_state[12]_net_1\, Y => N_151);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \rd_curr_state[1]\ : SLE
      port map(D => \rd_curr_state[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[1]_net_1\);
    
    \rd_curr_state_RNO[3]\ : CFG4
      generic map(INIT => x"080F")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, B => 
        AR_REQ_MI0, C => \rd_curr_state_ns_i_0[10]_net_1\, D => 
        N_149, Y => N_134_i);
    
    \AR_MASGNT_MI_xhdl1[1]\ : SLE
      port map(D => N_165_i, CLK => SDRCLK_c, EN => 
        \rd_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AR_MASGNT_IC(1));
    
    \AR_MASGNT_MI_xhdl1[0]\ : SLE
      port map(D => N_142_i, CLK => SDRCLK_c, EN => 
        \rd_curr_state_i[12]\, ALn => MSS_READY, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AR_MASGNT_IC(0));
    
    \AR_MASGNT_MI_xhdl1[3]\ : SLE
      port map(D => N_164_i, CLK => SDRCLK_c, EN => 
        \rd_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AR_MASGNT_IC(3));
    
    \rd_curr_state_ns_i_o2[10]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => \m0_lock_clear_read\, B => 
        \rd_curr_state[3]_net_1\, C => m0_rd_end, Y => N_149);
    
    \AR_MASGNT_MI_xhdl1_RNO[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \rd_curr_state[1]_net_1\, B => 
        \rd_curr_state[9]_net_1\, Y => N_163_i);
    
    \rd_curr_state_ns_a2_0[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \rd_curr_state[11]_net_1\, B => m0_rd_end, Y
         => N_158);
    
    \rd_curr_state_ns_i_0[10]\ : CFG4
      generic map(INIT => x"F0F1")

      port map(A => \rd_curr_state[3]_net_1\, B => 
        \rd_curr_state[13]_net_1\, C => N_158, D => N_151, Y => 
        \rd_curr_state_ns_i_0[10]_net_1\);
    
    \AR_MASGNT_MI_xhdl1[2]\ : SLE
      port map(D => N_163_i, CLK => SDRCLK_c, EN => 
        \rd_curr_state_i[12]\, ALn => MSS_READY, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => AR_MASGNT_IC(2));
    
    \rd_curr_state[10]\ : SLE
      port map(D => \rd_curr_state[10]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[10]_net_1\);
    
    m0_lock_clear_read : SLE
      port map(D => ARLOCK_MI0_i_0, CLK => SDRCLK_c, EN => 
        AR_REQ_MI0, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \m0_lock_clear_read\);
    
    \rd_curr_state_ns_a2[6]\ : CFG3
      generic map(INIT => x"08")

      port map(A => m0_rd_end, B => \rd_curr_state[11]_net_1\, C
         => AR_REQ_MI0, Y => \rd_curr_state_ns[6]\);
    
    \rd_curr_state[13]\ : SLE
      port map(D => \rd_curr_state_ns[0]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[13]_net_1\);
    
    \AR_MASGNT_MI_xhdl1_RNO[0]\ : CFG3
      generic map(INIT => x"31")

      port map(A => N_149, B => \rd_curr_state_ns[6]\, C => 
        \rd_curr_state[11]_net_1\, Y => N_142_i);
    
    \rd_curr_state[8]\ : SLE
      port map(D => \rd_curr_state[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[8]_net_1\);
    
    \rd_curr_state_ns[2]\ : CFG4
      generic map(INIT => x"F2F0")

      port map(A => AR_REQ_MI0, B => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, C => N_158, D => 
        N_152, Y => \rd_curr_state_ns[2]_net_1\);
    
    \rd_curr_state[9]\ : SLE
      port map(D => \rd_curr_state[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[9]_net_1\);
    
    \rd_curr_state[0]\ : SLE
      port map(D => \rd_curr_state[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rd_curr_state[0]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_rdmatrix_4Mto1S is

    port( ARSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1);
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARLOCK_MI0_i_0                       : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          ARBURST_MI0_0                        : in    std_logic;
          ARBURST_IS16_gated_0                 : out   std_logic;
          m0_rd_end                            : in    std_logic;
          ARVALID_MI0                          : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          ARVALID_IS16_gated                   : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_rdmatrix_4Mto1S;

architecture DEF_ARCH of axi_rdmatrix_4Mto1S is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component axi_RA_ARBITER
    port( AR_MASGNT_IC                         : out   std_logic_vector(3 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          ARLOCK_MI0_i_0                       : in    std_logic := 'U';
          m0_rd_end                            : in    std_logic := 'U';
          AR_REQ_MI0                           : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \ARBURST_IS_int[0]_net_1\, GND_net_1, 
        \ARSIZE_IS_int[0]_net_1\, \ARSIZE_IS_int[1]_net_1\, 
        \ARADDR_IS_int_xhdl14[22]_net_1\, arready_im0_int4, 
        \ARADDR_IS_int_xhdl14[23]_net_1\, 
        \ARADDR_IS_int_xhdl14[26]_net_1\, 
        \ARADDR_IS_int_xhdl14[27]_net_1\, \ARBURST_IS_int_3[0]\, 
        \ARSIZE_IS_int_3[0]\, \ARSIZE_IS_int_3[1]\, 
        \ARADDR_IS_int_xhdl14[7]_net_1\, 
        \ARADDR_IS_int_xhdl14[8]_net_1\, 
        \ARADDR_IS_int_xhdl14[9]_net_1\, 
        \ARADDR_IS_int_xhdl14[10]_net_1\, 
        \ARADDR_IS_int_xhdl14[11]_net_1\, 
        \ARADDR_IS_int_xhdl14[12]_net_1\, 
        \ARADDR_IS_int_xhdl14[13]_net_1\, 
        \ARADDR_IS_int_xhdl14[14]_net_1\, 
        \ARADDR_IS_int_xhdl14[15]_net_1\, 
        \ARADDR_IS_int_xhdl14[16]_net_1\, 
        \ARADDR_IS_int_xhdl14[17]_net_1\, 
        \ARADDR_IS_int_xhdl14[18]_net_1\, 
        \ARADDR_IS_int_xhdl14[19]_net_1\, 
        \ARADDR_IS_int_xhdl14[20]_net_1\, 
        \ARADDR_IS_int_xhdl14[21]_net_1\, 
        \ARADDR_IS_int_xhdl14[1]_net_1\, 
        \ARADDR_IS_int_xhdl14[2]_net_1\, 
        \ARADDR_IS_int_xhdl14[3]_net_1\, 
        \ARADDR_IS_int_xhdl14[4]_net_1\, 
        \ARADDR_IS_int_xhdl14[5]_net_1\, 
        \ARADDR_IS_int_xhdl14[6]_net_1\, \ARREADY_IM0_int\, 
        \ARVALID_IS_int\, ARVALID_IS_int_3, \AR_REQ_MI0\, 
        \AR_MASGNT_IC[3]\, \AR_MASGNT_IC[2]\, \AR_MASGNT_IC[1]\, 
        \AR_MASGNT_IC[0]\ : std_logic;

    for all : axi_RA_ARBITER
	Use entity work.axi_RA_ARBITER(DEF_ARCH);
begin 


    ARREADY_IM0_xhdl1 : SLE
      port map(D => \ARREADY_IM0_int\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ARREADY_IM0);
    
    \ARADDR_IS_xhdl6[16]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[16]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(16));
    
    \ARSIZE_IS_int[0]\ : SLE
      port map(D => \ARSIZE_IS_int_3[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARSIZE_IS_int[0]_net_1\);
    
    \ARADDR_IS_xhdl6[5]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[5]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(5));
    
    \ARADDR_IS_int_xhdl14[8]\ : SLE
      port map(D => ARADDR_MI0(8), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[8]_net_1\);
    
    \ARSIZE_IS_xhdl8[1]\ : SLE
      port map(D => \ARSIZE_IS_int[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ARSIZE_IS16_gated(1));
    
    \ARADDR_IS_xhdl6[26]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[26]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(26));
    
    \ARADDR_IS_xhdl6[9]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[9]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(9));
    
    \ARADDR_IS_xhdl6[8]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[8]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(8));
    
    \ARADDR_IS_int_xhdl14[26]\ : SLE
      port map(D => ARADDR_MI0(26), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[26]_net_1\);
    
    \ARADDR_IS_int_xhdl14[27]\ : SLE
      port map(D => ARADDR_MI0(27), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[27]_net_1\);
    
    \ARADDR_IS_int_xhdl14[20]\ : SLE
      port map(D => ARADDR_MI0(20), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[20]_net_1\);
    
    \ARADDR_IS_xhdl6[1]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[1]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(1));
    
    \ARADDR_IS_int_xhdl14[21]\ : SLE
      port map(D => ARADDR_MI0(21), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[21]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ARBURST_IS_xhdl9[0]\ : SLE
      port map(D => \ARBURST_IS_int[0]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ARBURST_IS16_gated_0);
    
    \ARADDR_IS_xhdl6[18]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[18]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(18));
    
    \ARADDR_IS_int_xhdl14[22]\ : SLE
      port map(D => ARADDR_MI0(22), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[22]_net_1\);
    
    \ARADDR_IS_int_xhdl14[9]\ : SLE
      port map(D => ARADDR_MI0(9), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[9]_net_1\);
    
    \ARADDR_IS_xhdl6[17]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[17]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(17));
    
    \ARADDR_IS_xhdl6[3]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[3]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(3));
    
    \ARADDR_IS_xhdl6[27]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[27]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(27));
    
    \ARADDR_IS_int_xhdl14[18]\ : SLE
      port map(D => ARADDR_MI0(18), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[18]_net_1\);
    
    \ARADDR_IS_int_xhdl14[2]\ : SLE
      port map(D => ARADDR_MI0(2), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[2]_net_1\);
    
    \ARSIZE_IS_int[1]\ : SLE
      port map(D => \ARSIZE_IS_int_3[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARSIZE_IS_int[1]_net_1\);
    
    ARVALID_IS_xhdl13 : SLE
      port map(D => \ARVALID_IS_int\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ARVALID_IS16_gated);
    
    \ARADDR_IS_xhdl6[10]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[10]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(10));
    
    \ARADDR_IS_int_xhdl14[4]\ : SLE
      port map(D => ARADDR_MI0(4), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[4]_net_1\);
    
    \ARADDR_IS_xhdl6[7]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[7]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(7));
    
    \ARADDR_IS_int_xhdl14[13]\ : SLE
      port map(D => ARADDR_MI0(13), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[13]_net_1\);
    
    \ARADDR_IS_xhdl6[20]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[20]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(20));
    
    \ARADDR_IS_int_xhdl14[15]\ : SLE
      port map(D => ARADDR_MI0(15), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[15]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \ARADDR_IS_xhdl6[2]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[2]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(2));
    
    \L1.ARVALID_IS_int_3\ : CFG2
      generic map(INIT => x"8")

      port map(A => arready_im0_int4, B => ARVALID_MI0, Y => 
        ARVALID_IS_int_3);
    
    \ARADDR_IS_int_xhdl14[7]\ : SLE
      port map(D => ARADDR_MI0(7), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[7]_net_1\);
    
    \L1.ARBURST_IS_int_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => arready_im0_int4, B => ARBURST_MI0_0, Y => 
        \ARBURST_IS_int_3[0]\);
    
    \ARADDR_IS_int_xhdl14[3]\ : SLE
      port map(D => ARADDR_MI0(3), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[3]_net_1\);
    
    \ARADDR_IS_int_xhdl14[14]\ : SLE
      port map(D => ARADDR_MI0(14), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[14]_net_1\);
    
    \L1.arready_im0_int4\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \AR_MASGNT_IC[3]\, B => \AR_MASGNT_IC[2]\, C
         => \AR_MASGNT_IC[1]\, D => \AR_MASGNT_IC[0]\, Y => 
        arready_im0_int4);
    
    URA_ARBITER0 : axi_RA_ARBITER
      port map(AR_MASGNT_IC(3) => \AR_MASGNT_IC[3]\, 
        AR_MASGNT_IC(2) => \AR_MASGNT_IC[2]\, AR_MASGNT_IC(1) => 
        \AR_MASGNT_IC[1]\, AR_MASGNT_IC(0) => \AR_MASGNT_IC[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, ARLOCK_MI0_i_0 => 
        ARLOCK_MI0_i_0, m0_rd_end => m0_rd_end, AR_REQ_MI0 => 
        \AR_REQ_MI0\, SDRCLK_c => SDRCLK_c, MSS_READY => 
        MSS_READY);
    
    \ARADDR_IS_int_xhdl14[16]\ : SLE
      port map(D => ARADDR_MI0(16), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[16]_net_1\);
    
    \ARADDR_IS_xhdl6[19]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[19]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(19));
    
    \ARSIZE_IS_xhdl8[0]\ : SLE
      port map(D => \ARSIZE_IS_int[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ARSIZE_IS16_gated(0));
    
    \ARADDR_IS_int_xhdl14[17]\ : SLE
      port map(D => ARADDR_MI0(17), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[17]_net_1\);
    
    \ARADDR_IS_int_xhdl14[10]\ : SLE
      port map(D => ARADDR_MI0(10), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[10]_net_1\);
    
    \ARADDR_IS_int_xhdl14[11]\ : SLE
      port map(D => ARADDR_MI0(11), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[11]_net_1\);
    
    \ARADDR_IS_int_xhdl14[19]\ : SLE
      port map(D => ARADDR_MI0(19), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[19]_net_1\);
    
    ARVALID_IS_int : SLE
      port map(D => ARVALID_IS_int_3, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARVALID_IS_int\);
    
    \ARADDR_IS_int_xhdl14[12]\ : SLE
      port map(D => ARADDR_MI0(12), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[12]_net_1\);
    
    AR_REQ_MI0 : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_ARVALID, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AR_REQ_MI0\);
    
    \ARADDR_IS_xhdl6[13]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[13]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(13));
    
    \ARADDR_IS_xhdl6[6]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[6]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(6));
    
    \ARADDR_IS_xhdl6[15]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[15]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(15));
    
    \L1.ARSIZE_IS_int_3[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => arready_im0_int4, B => ARSIZE_MI0(1), Y => 
        \ARSIZE_IS_int_3[1]\);
    
    \ARADDR_IS_xhdl6[4]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[4]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(4));
    
    \ARADDR_IS_xhdl6[23]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[23]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(23));
    
    \ARADDR_IS_xhdl6[14]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[14]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(14));
    
    \ARADDR_IS_xhdl6[12]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[12]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(12));
    
    \ARBURST_IS_int[0]\ : SLE
      port map(D => \ARBURST_IS_int_3[0]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARBURST_IS_int[0]_net_1\);
    
    \ARADDR_IS_xhdl6[22]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[22]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(22));
    
    ARREADY_IM0_int : CFG3
      generic map(INIT => x"80")

      port map(A => COREAXI_0_AXImslave16_ARVALID, B => 
        arready_im0_int4, C => COREAXI_0_AXImslave16_ARREADY, Y
         => \ARREADY_IM0_int\);
    
    \ARADDR_IS_int_xhdl14[23]\ : SLE
      port map(D => ARADDR_MI0(23), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[23]_net_1\);
    
    \ARADDR_IS_int_xhdl14[1]\ : SLE
      port map(D => ARADDR_MI0(1), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[1]_net_1\);
    
    \ARADDR_IS_xhdl6[11]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[11]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(11));
    
    \L1.ARSIZE_IS_int_3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => arready_im0_int4, B => ARSIZE_MI0(0), Y => 
        \ARSIZE_IS_int_3[0]\);
    
    \ARADDR_IS_int_xhdl14[6]\ : SLE
      port map(D => ARADDR_MI0(6), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[6]_net_1\);
    
    \ARADDR_IS_xhdl6[21]\ : SLE
      port map(D => \ARADDR_IS_int_xhdl14[21]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ARADDR_IS16_gated(21));
    
    \ARADDR_IS_int_xhdl14[5]\ : SLE
      port map(D => ARADDR_MI0(5), CLK => SDRCLK_c, EN => 
        arready_im0_int4, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS_int_xhdl14[5]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_ra_channel is

    port( ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1);
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          ARBURST_IS16_gated_0                 : out   std_logic;
          ARBURST_MI0_0                        : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          ARLOCK_MI0_i_0                       : in    std_logic;
          MSS_READY                            : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          ARREADY_IM0                          : out   std_logic;
          ARVALID_IS16_gated                   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic;
          ARVALID_MI0                          : in    std_logic;
          m0_rd_end                            : in    std_logic
        );

end axi_ra_channel;

architecture DEF_ARCH of axi_ra_channel is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component axi_rdmatrix_4Mto1S
    port( ARSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARLOCK_MI0_i_0                       : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          ARBURST_MI0_0                        : in    std_logic := 'U';
          ARBURST_IS16_gated_0                 : out   std_logic;
          m0_rd_end                            : in    std_logic := 'U';
          ARVALID_MI0                          : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          ARVALID_IS16_gated                   : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : axi_rdmatrix_4Mto1S
	Use entity work.axi_rdmatrix_4Mto1S(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \L1.inst_rdmatrix_4Mto1S\ : axi_rdmatrix_4Mto1S
      port map(ARSIZE_MI0(1) => ARSIZE_MI0(1), ARSIZE_MI0(0) => 
        ARSIZE_MI0(0), ARADDR_IS16_gated(27) => 
        ARADDR_IS16_gated(27), ARADDR_IS16_gated(26) => 
        ARADDR_IS16_gated(26), ARADDR_IS16_gated(25) => nc2, 
        ARADDR_IS16_gated(24) => nc4, ARADDR_IS16_gated(23) => 
        ARADDR_IS16_gated(23), ARADDR_IS16_gated(22) => 
        ARADDR_IS16_gated(22), ARADDR_IS16_gated(21) => 
        ARADDR_IS16_gated(21), ARADDR_IS16_gated(20) => 
        ARADDR_IS16_gated(20), ARADDR_IS16_gated(19) => 
        ARADDR_IS16_gated(19), ARADDR_IS16_gated(18) => 
        ARADDR_IS16_gated(18), ARADDR_IS16_gated(17) => 
        ARADDR_IS16_gated(17), ARADDR_IS16_gated(16) => 
        ARADDR_IS16_gated(16), ARADDR_IS16_gated(15) => 
        ARADDR_IS16_gated(15), ARADDR_IS16_gated(14) => 
        ARADDR_IS16_gated(14), ARADDR_IS16_gated(13) => 
        ARADDR_IS16_gated(13), ARADDR_IS16_gated(12) => 
        ARADDR_IS16_gated(12), ARADDR_IS16_gated(11) => 
        ARADDR_IS16_gated(11), ARADDR_IS16_gated(10) => 
        ARADDR_IS16_gated(10), ARADDR_IS16_gated(9) => 
        ARADDR_IS16_gated(9), ARADDR_IS16_gated(8) => 
        ARADDR_IS16_gated(8), ARADDR_IS16_gated(7) => 
        ARADDR_IS16_gated(7), ARADDR_IS16_gated(6) => 
        ARADDR_IS16_gated(6), ARADDR_IS16_gated(5) => 
        ARADDR_IS16_gated(5), ARADDR_IS16_gated(4) => 
        ARADDR_IS16_gated(4), ARADDR_IS16_gated(3) => 
        ARADDR_IS16_gated(3), ARADDR_IS16_gated(2) => 
        ARADDR_IS16_gated(2), ARADDR_IS16_gated(1) => 
        ARADDR_IS16_gated(1), ARADDR_MI0(27) => ARADDR_MI0(27), 
        ARADDR_MI0(26) => ARADDR_MI0(26), ARADDR_MI0(25) => nc3, 
        ARADDR_MI0(24) => nc1, ARADDR_MI0(23) => ARADDR_MI0(23), 
        ARADDR_MI0(22) => ARADDR_MI0(22), ARADDR_MI0(21) => 
        ARADDR_MI0(21), ARADDR_MI0(20) => ARADDR_MI0(20), 
        ARADDR_MI0(19) => ARADDR_MI0(19), ARADDR_MI0(18) => 
        ARADDR_MI0(18), ARADDR_MI0(17) => ARADDR_MI0(17), 
        ARADDR_MI0(16) => ARADDR_MI0(16), ARADDR_MI0(15) => 
        ARADDR_MI0(15), ARADDR_MI0(14) => ARADDR_MI0(14), 
        ARADDR_MI0(13) => ARADDR_MI0(13), ARADDR_MI0(12) => 
        ARADDR_MI0(12), ARADDR_MI0(11) => ARADDR_MI0(11), 
        ARADDR_MI0(10) => ARADDR_MI0(10), ARADDR_MI0(9) => 
        ARADDR_MI0(9), ARADDR_MI0(8) => ARADDR_MI0(8), 
        ARADDR_MI0(7) => ARADDR_MI0(7), ARADDR_MI0(6) => 
        ARADDR_MI0(6), ARADDR_MI0(5) => ARADDR_MI0(5), 
        ARADDR_MI0(4) => ARADDR_MI0(4), ARADDR_MI0(3) => 
        ARADDR_MI0(3), ARADDR_MI0(2) => ARADDR_MI0(2), 
        ARADDR_MI0(1) => ARADDR_MI0(1), ARSIZE_IS16_gated(1) => 
        ARSIZE_IS16_gated(1), ARSIZE_IS16_gated(0) => 
        ARSIZE_IS16_gated(0), ARLOCK_MI0_i_0 => ARLOCK_MI0_i_0, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, ARBURST_MI0_0 => 
        ARBURST_MI0_0, ARBURST_IS16_gated_0 => 
        ARBURST_IS16_gated_0, m0_rd_end => m0_rd_end, ARVALID_MI0
         => ARVALID_MI0, COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, 
        COREAXI_0_AXImslave16_ARVALID => 
        COREAXI_0_AXImslave16_ARVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, ARVALID_IS16_gated
         => ARVALID_IS16_gated, ARREADY_IM0 => ARREADY_IM0, 
        SDRCLK_c => SDRCLK_c, MSS_READY => MSS_READY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_matrix_s is

    port( ARSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1);
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          WSTRB_IS16_gated                     : out   std_logic_vector(7 downto 0);
          WDATA_IS16_gated                     : out   std_logic_vector(63 downto 0);
          WSTRB_MI0                            : in    std_logic_vector(7 downto 0);
          WDATA_MI0                            : in    std_logic_vector(63 downto 0);
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1);
          AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARLOCK_MI0_i_0                       : in    std_logic;
          ARBURST_MI0_0                        : in    std_logic;
          ARBURST_IS16_gated_0                 : out   std_logic;
          AWLOCK_MI0_i_0                       : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          m0_rd_end                            : in    std_logic;
          ARVALID_MI0                          : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          ARVALID_IS16_gated                   : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          WREADY_IM0                           : out   std_logic;
          WVALID_IS16_gated                    : out   std_logic;
          WVALID_MI0                           : in    std_logic;
          WREADY_SI16                          : in    std_logic;
          m0_wr_end                            : in    std_logic;
          AWREADY_SI16                         : in    std_logic;
          AWVALID_MI0                          : in    std_logic;
          N_75_i                               : in    std_logic;
          AWVALID_IS16_gated                   : out   std_logic;
          AWREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_matrix_s;

architecture DEF_ARCH of axi_matrix_s is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component axi_wa_channel
    port( AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          MST_WRGNT_NUM_0                      : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          AWLOCK_MI0_i_0                       : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          AWREADY_IM0                          : out   std_logic;
          AWVALID_IS16_gated                   : out   std_logic;
          N_75_i                               : in    std_logic := 'U';
          AWVALID_MI0                          : in    std_logic := 'U';
          AWREADY_SI16                         : in    std_logic := 'U';
          m0_wr_end                            : in    std_logic := 'U'
        );
  end component;

  component axi_wd_channel
    port( WDATA_MI0         : in    std_logic_vector(63 downto 0) := (others => 'U');
          WSTRB_MI0         : in    std_logic_vector(7 downto 0) := (others => 'U');
          WDATA_IS16_gated  : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated  : out   std_logic_vector(7 downto 0);
          MST_WRGNT_NUM_0   : in    std_logic := 'U';
          WREADY_SI16       : in    std_logic := 'U';
          WVALID_MI0        : in    std_logic := 'U';
          WVALID_IS16_gated : out   std_logic;
          WREADY_IM0        : out   std_logic;
          SDRCLK_c          : in    std_logic := 'U';
          MSS_READY         : in    std_logic := 'U'
        );
  end component;

  component axi_ra_channel
    port( ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          ARBURST_IS16_gated_0                 : out   std_logic;
          ARBURST_MI0_0                        : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          ARLOCK_MI0_i_0                       : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          ARREADY_IM0                          : out   std_logic;
          ARVALID_IS16_gated                   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic := 'U';
          ARVALID_MI0                          : in    std_logic := 'U';
          m0_rd_end                            : in    std_logic := 'U'
        );
  end component;

    signal \MST_WRGNT_NUM[0]\, GND_net_1, VCC_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

    for all : axi_wa_channel
	Use entity work.axi_wa_channel(DEF_ARCH);
    for all : axi_wd_channel
	Use entity work.axi_wd_channel(DEF_ARCH);
    for all : axi_ra_channel
	Use entity work.axi_ra_channel(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    inst_wa_channel : axi_wa_channel
      port map(AWSIZE_IS16_gated(1) => AWSIZE_IS16_gated(1), 
        AWSIZE_IS16_gated(0) => AWSIZE_IS16_gated(0), 
        AWADDR_MI0(27) => AWADDR_MI0(27), AWADDR_MI0(26) => 
        AWADDR_MI0(26), AWADDR_MI0(25) => nc8, AWADDR_MI0(24) => 
        nc7, AWADDR_MI0(23) => AWADDR_MI0(23), AWADDR_MI0(22) => 
        AWADDR_MI0(22), AWADDR_MI0(21) => AWADDR_MI0(21), 
        AWADDR_MI0(20) => AWADDR_MI0(20), AWADDR_MI0(19) => 
        AWADDR_MI0(19), AWADDR_MI0(18) => AWADDR_MI0(18), 
        AWADDR_MI0(17) => AWADDR_MI0(17), AWADDR_MI0(16) => 
        AWADDR_MI0(16), AWADDR_MI0(15) => AWADDR_MI0(15), 
        AWADDR_MI0(14) => AWADDR_MI0(14), AWADDR_MI0(13) => 
        AWADDR_MI0(13), AWADDR_MI0(12) => AWADDR_MI0(12), 
        AWADDR_MI0(11) => AWADDR_MI0(11), AWADDR_MI0(10) => 
        AWADDR_MI0(10), AWADDR_MI0(9) => AWADDR_MI0(9), 
        AWADDR_MI0(8) => AWADDR_MI0(8), AWADDR_MI0(7) => 
        AWADDR_MI0(7), AWADDR_MI0(6) => AWADDR_MI0(6), 
        AWADDR_MI0(5) => AWADDR_MI0(5), AWADDR_MI0(4) => 
        AWADDR_MI0(4), AWADDR_MI0(3) => AWADDR_MI0(3), 
        AWADDR_MI0(2) => AWADDR_MI0(2), AWADDR_MI0(1) => 
        AWADDR_MI0(1), AWADDR_IS16_gated(27) => 
        AWADDR_IS16_gated(27), AWADDR_IS16_gated(26) => 
        AWADDR_IS16_gated(26), AWADDR_IS16_gated(25) => nc6, 
        AWADDR_IS16_gated(24) => nc2, AWADDR_IS16_gated(23) => 
        AWADDR_IS16_gated(23), AWADDR_IS16_gated(22) => 
        AWADDR_IS16_gated(22), AWADDR_IS16_gated(21) => 
        AWADDR_IS16_gated(21), AWADDR_IS16_gated(20) => 
        AWADDR_IS16_gated(20), AWADDR_IS16_gated(19) => 
        AWADDR_IS16_gated(19), AWADDR_IS16_gated(18) => 
        AWADDR_IS16_gated(18), AWADDR_IS16_gated(17) => 
        AWADDR_IS16_gated(17), AWADDR_IS16_gated(16) => 
        AWADDR_IS16_gated(16), AWADDR_IS16_gated(15) => 
        AWADDR_IS16_gated(15), AWADDR_IS16_gated(14) => 
        AWADDR_IS16_gated(14), AWADDR_IS16_gated(13) => 
        AWADDR_IS16_gated(13), AWADDR_IS16_gated(12) => 
        AWADDR_IS16_gated(12), AWADDR_IS16_gated(11) => 
        AWADDR_IS16_gated(11), AWADDR_IS16_gated(10) => 
        AWADDR_IS16_gated(10), AWADDR_IS16_gated(9) => 
        AWADDR_IS16_gated(9), AWADDR_IS16_gated(8) => 
        AWADDR_IS16_gated(8), AWADDR_IS16_gated(7) => 
        AWADDR_IS16_gated(7), AWADDR_IS16_gated(6) => 
        AWADDR_IS16_gated(6), AWADDR_IS16_gated(5) => 
        AWADDR_IS16_gated(5), AWADDR_IS16_gated(4) => 
        AWADDR_IS16_gated(4), AWADDR_IS16_gated(3) => 
        AWADDR_IS16_gated(3), AWADDR_IS16_gated(2) => 
        AWADDR_IS16_gated(2), AWADDR_IS16_gated(1) => 
        AWADDR_IS16_gated(1), AWSIZE_MI0(1) => AWSIZE_MI0(1), 
        AWSIZE_MI0(0) => AWSIZE_MI0(0), MST_WRGNT_NUM_0 => 
        \MST_WRGNT_NUM[0]\, COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0
         => COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, AWLOCK_MI0_i_0
         => AWLOCK_MI0_i_0, MSS_READY => MSS_READY, SDRCLK_c => 
        SDRCLK_c, AWREADY_IM0 => AWREADY_IM0, AWVALID_IS16_gated
         => AWVALID_IS16_gated, N_75_i => N_75_i, AWVALID_MI0 => 
        AWVALID_MI0, AWREADY_SI16 => AWREADY_SI16, m0_wr_end => 
        m0_wr_end);
    
    inst_wd_channel : axi_wd_channel
      port map(WDATA_MI0(63) => WDATA_MI0(63), WDATA_MI0(62) => 
        WDATA_MI0(62), WDATA_MI0(61) => WDATA_MI0(61), 
        WDATA_MI0(60) => WDATA_MI0(60), WDATA_MI0(59) => 
        WDATA_MI0(59), WDATA_MI0(58) => WDATA_MI0(58), 
        WDATA_MI0(57) => WDATA_MI0(57), WDATA_MI0(56) => 
        WDATA_MI0(56), WDATA_MI0(55) => WDATA_MI0(55), 
        WDATA_MI0(54) => WDATA_MI0(54), WDATA_MI0(53) => 
        WDATA_MI0(53), WDATA_MI0(52) => WDATA_MI0(52), 
        WDATA_MI0(51) => WDATA_MI0(51), WDATA_MI0(50) => 
        WDATA_MI0(50), WDATA_MI0(49) => WDATA_MI0(49), 
        WDATA_MI0(48) => WDATA_MI0(48), WDATA_MI0(47) => 
        WDATA_MI0(47), WDATA_MI0(46) => WDATA_MI0(46), 
        WDATA_MI0(45) => WDATA_MI0(45), WDATA_MI0(44) => 
        WDATA_MI0(44), WDATA_MI0(43) => WDATA_MI0(43), 
        WDATA_MI0(42) => WDATA_MI0(42), WDATA_MI0(41) => 
        WDATA_MI0(41), WDATA_MI0(40) => WDATA_MI0(40), 
        WDATA_MI0(39) => WDATA_MI0(39), WDATA_MI0(38) => 
        WDATA_MI0(38), WDATA_MI0(37) => WDATA_MI0(37), 
        WDATA_MI0(36) => WDATA_MI0(36), WDATA_MI0(35) => 
        WDATA_MI0(35), WDATA_MI0(34) => WDATA_MI0(34), 
        WDATA_MI0(33) => WDATA_MI0(33), WDATA_MI0(32) => 
        WDATA_MI0(32), WDATA_MI0(31) => WDATA_MI0(31), 
        WDATA_MI0(30) => WDATA_MI0(30), WDATA_MI0(29) => 
        WDATA_MI0(29), WDATA_MI0(28) => WDATA_MI0(28), 
        WDATA_MI0(27) => WDATA_MI0(27), WDATA_MI0(26) => 
        WDATA_MI0(26), WDATA_MI0(25) => WDATA_MI0(25), 
        WDATA_MI0(24) => WDATA_MI0(24), WDATA_MI0(23) => 
        WDATA_MI0(23), WDATA_MI0(22) => WDATA_MI0(22), 
        WDATA_MI0(21) => WDATA_MI0(21), WDATA_MI0(20) => 
        WDATA_MI0(20), WDATA_MI0(19) => WDATA_MI0(19), 
        WDATA_MI0(18) => WDATA_MI0(18), WDATA_MI0(17) => 
        WDATA_MI0(17), WDATA_MI0(16) => WDATA_MI0(16), 
        WDATA_MI0(15) => WDATA_MI0(15), WDATA_MI0(14) => 
        WDATA_MI0(14), WDATA_MI0(13) => WDATA_MI0(13), 
        WDATA_MI0(12) => WDATA_MI0(12), WDATA_MI0(11) => 
        WDATA_MI0(11), WDATA_MI0(10) => WDATA_MI0(10), 
        WDATA_MI0(9) => WDATA_MI0(9), WDATA_MI0(8) => 
        WDATA_MI0(8), WDATA_MI0(7) => WDATA_MI0(7), WDATA_MI0(6)
         => WDATA_MI0(6), WDATA_MI0(5) => WDATA_MI0(5), 
        WDATA_MI0(4) => WDATA_MI0(4), WDATA_MI0(3) => 
        WDATA_MI0(3), WDATA_MI0(2) => WDATA_MI0(2), WDATA_MI0(1)
         => WDATA_MI0(1), WDATA_MI0(0) => WDATA_MI0(0), 
        WSTRB_MI0(7) => WSTRB_MI0(7), WSTRB_MI0(6) => 
        WSTRB_MI0(6), WSTRB_MI0(5) => WSTRB_MI0(5), WSTRB_MI0(4)
         => WSTRB_MI0(4), WSTRB_MI0(3) => WSTRB_MI0(3), 
        WSTRB_MI0(2) => WSTRB_MI0(2), WSTRB_MI0(1) => 
        WSTRB_MI0(1), WSTRB_MI0(0) => WSTRB_MI0(0), 
        WDATA_IS16_gated(63) => WDATA_IS16_gated(63), 
        WDATA_IS16_gated(62) => WDATA_IS16_gated(62), 
        WDATA_IS16_gated(61) => WDATA_IS16_gated(61), 
        WDATA_IS16_gated(60) => WDATA_IS16_gated(60), 
        WDATA_IS16_gated(59) => WDATA_IS16_gated(59), 
        WDATA_IS16_gated(58) => WDATA_IS16_gated(58), 
        WDATA_IS16_gated(57) => WDATA_IS16_gated(57), 
        WDATA_IS16_gated(56) => WDATA_IS16_gated(56), 
        WDATA_IS16_gated(55) => WDATA_IS16_gated(55), 
        WDATA_IS16_gated(54) => WDATA_IS16_gated(54), 
        WDATA_IS16_gated(53) => WDATA_IS16_gated(53), 
        WDATA_IS16_gated(52) => WDATA_IS16_gated(52), 
        WDATA_IS16_gated(51) => WDATA_IS16_gated(51), 
        WDATA_IS16_gated(50) => WDATA_IS16_gated(50), 
        WDATA_IS16_gated(49) => WDATA_IS16_gated(49), 
        WDATA_IS16_gated(48) => WDATA_IS16_gated(48), 
        WDATA_IS16_gated(47) => WDATA_IS16_gated(47), 
        WDATA_IS16_gated(46) => WDATA_IS16_gated(46), 
        WDATA_IS16_gated(45) => WDATA_IS16_gated(45), 
        WDATA_IS16_gated(44) => WDATA_IS16_gated(44), 
        WDATA_IS16_gated(43) => WDATA_IS16_gated(43), 
        WDATA_IS16_gated(42) => WDATA_IS16_gated(42), 
        WDATA_IS16_gated(41) => WDATA_IS16_gated(41), 
        WDATA_IS16_gated(40) => WDATA_IS16_gated(40), 
        WDATA_IS16_gated(39) => WDATA_IS16_gated(39), 
        WDATA_IS16_gated(38) => WDATA_IS16_gated(38), 
        WDATA_IS16_gated(37) => WDATA_IS16_gated(37), 
        WDATA_IS16_gated(36) => WDATA_IS16_gated(36), 
        WDATA_IS16_gated(35) => WDATA_IS16_gated(35), 
        WDATA_IS16_gated(34) => WDATA_IS16_gated(34), 
        WDATA_IS16_gated(33) => WDATA_IS16_gated(33), 
        WDATA_IS16_gated(32) => WDATA_IS16_gated(32), 
        WDATA_IS16_gated(31) => WDATA_IS16_gated(31), 
        WDATA_IS16_gated(30) => WDATA_IS16_gated(30), 
        WDATA_IS16_gated(29) => WDATA_IS16_gated(29), 
        WDATA_IS16_gated(28) => WDATA_IS16_gated(28), 
        WDATA_IS16_gated(27) => WDATA_IS16_gated(27), 
        WDATA_IS16_gated(26) => WDATA_IS16_gated(26), 
        WDATA_IS16_gated(25) => WDATA_IS16_gated(25), 
        WDATA_IS16_gated(24) => WDATA_IS16_gated(24), 
        WDATA_IS16_gated(23) => WDATA_IS16_gated(23), 
        WDATA_IS16_gated(22) => WDATA_IS16_gated(22), 
        WDATA_IS16_gated(21) => WDATA_IS16_gated(21), 
        WDATA_IS16_gated(20) => WDATA_IS16_gated(20), 
        WDATA_IS16_gated(19) => WDATA_IS16_gated(19), 
        WDATA_IS16_gated(18) => WDATA_IS16_gated(18), 
        WDATA_IS16_gated(17) => WDATA_IS16_gated(17), 
        WDATA_IS16_gated(16) => WDATA_IS16_gated(16), 
        WDATA_IS16_gated(15) => WDATA_IS16_gated(15), 
        WDATA_IS16_gated(14) => WDATA_IS16_gated(14), 
        WDATA_IS16_gated(13) => WDATA_IS16_gated(13), 
        WDATA_IS16_gated(12) => WDATA_IS16_gated(12), 
        WDATA_IS16_gated(11) => WDATA_IS16_gated(11), 
        WDATA_IS16_gated(10) => WDATA_IS16_gated(10), 
        WDATA_IS16_gated(9) => WDATA_IS16_gated(9), 
        WDATA_IS16_gated(8) => WDATA_IS16_gated(8), 
        WDATA_IS16_gated(7) => WDATA_IS16_gated(7), 
        WDATA_IS16_gated(6) => WDATA_IS16_gated(6), 
        WDATA_IS16_gated(5) => WDATA_IS16_gated(5), 
        WDATA_IS16_gated(4) => WDATA_IS16_gated(4), 
        WDATA_IS16_gated(3) => WDATA_IS16_gated(3), 
        WDATA_IS16_gated(2) => WDATA_IS16_gated(2), 
        WDATA_IS16_gated(1) => WDATA_IS16_gated(1), 
        WDATA_IS16_gated(0) => WDATA_IS16_gated(0), 
        WSTRB_IS16_gated(7) => WSTRB_IS16_gated(7), 
        WSTRB_IS16_gated(6) => WSTRB_IS16_gated(6), 
        WSTRB_IS16_gated(5) => WSTRB_IS16_gated(5), 
        WSTRB_IS16_gated(4) => WSTRB_IS16_gated(4), 
        WSTRB_IS16_gated(3) => WSTRB_IS16_gated(3), 
        WSTRB_IS16_gated(2) => WSTRB_IS16_gated(2), 
        WSTRB_IS16_gated(1) => WSTRB_IS16_gated(1), 
        WSTRB_IS16_gated(0) => WSTRB_IS16_gated(0), 
        MST_WRGNT_NUM_0 => \MST_WRGNT_NUM[0]\, WREADY_SI16 => 
        WREADY_SI16, WVALID_MI0 => WVALID_MI0, WVALID_IS16_gated
         => WVALID_IS16_gated, WREADY_IM0 => WREADY_IM0, SDRCLK_c
         => SDRCLK_c, MSS_READY => MSS_READY);
    
    inst_ra_channel : axi_ra_channel
      port map(ARSIZE_IS16_gated(1) => ARSIZE_IS16_gated(1), 
        ARSIZE_IS16_gated(0) => ARSIZE_IS16_gated(0), 
        ARADDR_MI0(27) => ARADDR_MI0(27), ARADDR_MI0(26) => 
        ARADDR_MI0(26), ARADDR_MI0(25) => nc5, ARADDR_MI0(24) => 
        nc4, ARADDR_MI0(23) => ARADDR_MI0(23), ARADDR_MI0(22) => 
        ARADDR_MI0(22), ARADDR_MI0(21) => ARADDR_MI0(21), 
        ARADDR_MI0(20) => ARADDR_MI0(20), ARADDR_MI0(19) => 
        ARADDR_MI0(19), ARADDR_MI0(18) => ARADDR_MI0(18), 
        ARADDR_MI0(17) => ARADDR_MI0(17), ARADDR_MI0(16) => 
        ARADDR_MI0(16), ARADDR_MI0(15) => ARADDR_MI0(15), 
        ARADDR_MI0(14) => ARADDR_MI0(14), ARADDR_MI0(13) => 
        ARADDR_MI0(13), ARADDR_MI0(12) => ARADDR_MI0(12), 
        ARADDR_MI0(11) => ARADDR_MI0(11), ARADDR_MI0(10) => 
        ARADDR_MI0(10), ARADDR_MI0(9) => ARADDR_MI0(9), 
        ARADDR_MI0(8) => ARADDR_MI0(8), ARADDR_MI0(7) => 
        ARADDR_MI0(7), ARADDR_MI0(6) => ARADDR_MI0(6), 
        ARADDR_MI0(5) => ARADDR_MI0(5), ARADDR_MI0(4) => 
        ARADDR_MI0(4), ARADDR_MI0(3) => ARADDR_MI0(3), 
        ARADDR_MI0(2) => ARADDR_MI0(2), ARADDR_MI0(1) => 
        ARADDR_MI0(1), ARADDR_IS16_gated(27) => 
        ARADDR_IS16_gated(27), ARADDR_IS16_gated(26) => 
        ARADDR_IS16_gated(26), ARADDR_IS16_gated(25) => nc3, 
        ARADDR_IS16_gated(24) => nc1, ARADDR_IS16_gated(23) => 
        ARADDR_IS16_gated(23), ARADDR_IS16_gated(22) => 
        ARADDR_IS16_gated(22), ARADDR_IS16_gated(21) => 
        ARADDR_IS16_gated(21), ARADDR_IS16_gated(20) => 
        ARADDR_IS16_gated(20), ARADDR_IS16_gated(19) => 
        ARADDR_IS16_gated(19), ARADDR_IS16_gated(18) => 
        ARADDR_IS16_gated(18), ARADDR_IS16_gated(17) => 
        ARADDR_IS16_gated(17), ARADDR_IS16_gated(16) => 
        ARADDR_IS16_gated(16), ARADDR_IS16_gated(15) => 
        ARADDR_IS16_gated(15), ARADDR_IS16_gated(14) => 
        ARADDR_IS16_gated(14), ARADDR_IS16_gated(13) => 
        ARADDR_IS16_gated(13), ARADDR_IS16_gated(12) => 
        ARADDR_IS16_gated(12), ARADDR_IS16_gated(11) => 
        ARADDR_IS16_gated(11), ARADDR_IS16_gated(10) => 
        ARADDR_IS16_gated(10), ARADDR_IS16_gated(9) => 
        ARADDR_IS16_gated(9), ARADDR_IS16_gated(8) => 
        ARADDR_IS16_gated(8), ARADDR_IS16_gated(7) => 
        ARADDR_IS16_gated(7), ARADDR_IS16_gated(6) => 
        ARADDR_IS16_gated(6), ARADDR_IS16_gated(5) => 
        ARADDR_IS16_gated(5), ARADDR_IS16_gated(4) => 
        ARADDR_IS16_gated(4), ARADDR_IS16_gated(3) => 
        ARADDR_IS16_gated(3), ARADDR_IS16_gated(2) => 
        ARADDR_IS16_gated(2), ARADDR_IS16_gated(1) => 
        ARADDR_IS16_gated(1), ARSIZE_MI0(1) => ARSIZE_MI0(1), 
        ARSIZE_MI0(0) => ARSIZE_MI0(0), ARBURST_IS16_gated_0 => 
        ARBURST_IS16_gated_0, ARBURST_MI0_0 => ARBURST_MI0_0, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, ARLOCK_MI0_i_0 => 
        ARLOCK_MI0_i_0, MSS_READY => MSS_READY, SDRCLK_c => 
        SDRCLK_c, ARREADY_IM0 => ARREADY_IM0, ARVALID_IS16_gated
         => ARVALID_IS16_gated, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, 
        COREAXI_0_AXImslave16_ARVALID => 
        COREAXI_0_AXImslave16_ARVALID, 
        COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, ARVALID_MI0 => ARVALID_MI0, 
        m0_rd_end => m0_rd_end);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_rdmatrix_16Sto1M is

    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          axi_state_0                        : in    std_logic;
          RDATA_reg_3                        : in    std_logic;
          RDATA_reg_0                        : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic;
          N_3297                             : in    std_logic;
          RREADY_MI0                         : in    std_logic;
          N_389                              : in    std_logic;
          N_74                               : in    std_logic;
          N_3167_i                           : out   std_logic;
          N_23                               : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic;
          RVALID_IM0                         : out   std_logic;
          RLAST_IM0                          : out   std_logic;
          N_3170_i                           : in    std_logic;
          N_39                               : in    std_logic;
          N_78_mux_i                         : in    std_logic;
          N_79_mux_i                         : in    std_logic;
          N_80_mux_i                         : in    std_logic;
          N_70_mux_i                         : in    std_logic;
          N_71_mux_i                         : in    std_logic;
          N_72_mux_i                         : in    std_logic;
          N_3094_i                           : in    std_logic;
          N_3096_i                           : in    std_logic;
          N_3098_i                           : in    std_logic;
          N_3100_i                           : in    std_logic;
          N_3102_i                           : in    std_logic;
          N_3169_i                           : in    std_logic;
          N_3066_i                           : in    std_logic;
          N_67_mux_i                         : in    std_logic;
          N_68_mux_i                         : in    std_logic;
          N_69_mux_i                         : in    std_logic;
          N_75_mux_i                         : in    std_logic;
          N_76_mux_i                         : in    std_logic;
          N_77_mux_i                         : in    std_logic;
          i22_mux_2_i                        : in    std_logic;
          i22_mux_3_i                        : in    std_logic;
          i22_mux_4_i                        : in    std_logic;
          i22_mux_5_i                        : in    std_logic;
          N_8_i                              : in    std_logic;
          i17_mux_2_i                        : in    std_logic;
          N_3064_i                           : in    std_logic;
          N_3092_i                           : in    std_logic;
          i17_mux_i                          : in    std_logic;
          i17_mux_0_i                        : in    std_logic;
          i17_mux_1_i                        : in    std_logic;
          i22_mux_i                          : in    std_logic;
          i22_mux_0_i                        : in    std_logic;
          i22_mux_1_i                        : in    std_logic;
          SDRCLK_c                           : in    std_logic;
          MSS_READY                          : in    std_logic
        );

end axi_rdmatrix_16Sto1M;

architecture DEF_ARCH of axi_rdmatrix_16Sto1M is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1, 
        \COREAXI_0_AXImslave16_RDATA_m[43]\, 
        \COREAXI_0_AXImslave16_RDATA_m[46]\, 
        \curr_state[5]_net_1\, N_391_i, \curr_state[0]_net_1\, 
        N_384_i, COREAXI_0_AXImslave16_RLAST_m, \RVALID_IM0\, 
        rvalid_im_int_xhdl42_1, \RVALID_IM_r\, \N_3167_i\, N_3163
         : std_logic;

begin 

    N_3167_i <= \N_3167_i\;
    RVALID_IM0 <= \RVALID_IM0\;

    \curr_state_ns_i_0_o2[5]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_389, B => axi_state_0, Y => N_3163);
    
    \curr_state_RNO[5]\ : CFG4
      generic map(INIT => x"E2C0")

      port map(A => \RVALID_IM_r\, B => \curr_state[5]_net_1\, C
         => N_3163, D => RREADY_MI0, Y => N_391_i);
    
    RREADY_IS16_i_i_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => \RVALID_IM_r\, B => \curr_state[0]_net_1\, C
         => COREAHBLTOAXI_0_AXIMasterIF_RREADY, D => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, Y => N_23);
    
    \RDATA_IM_xhdl4[58]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_58, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(58));
    
    \RDATA_IM_xhdl4[30]\ : SLE
      port map(D => N_68_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(30));
    
    \RDATA_IM_xhdl4[61]\ : SLE
      port map(D => i17_mux_1_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(61));
    
    \RDATA_IM_xhdl4[5]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_5, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(5));
    
    \RDATA_IM_xhdl4[8]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_8, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(8));
    
    \RDATA_IM_xhdl4[40]\ : SLE
      port map(D => N_3094_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(40));
    
    \RDATA_IM_xhdl4[26]\ : SLE
      port map(D => N_77_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(26));
    
    \RDATA_IM_xhdl4[22]\ : SLE
      port map(D => N_80_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(22));
    
    \RDATA_IM_xhdl4[16]\ : SLE
      port map(D => N_72_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(16));
    
    \RDATA_IM_xhdl4[12]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_12, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(12));
    
    \RDATA_IM_xhdl4[59]\ : SLE
      port map(D => i22_mux_0_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(59));
    
    \RDATA_IM_xhdl4[57]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_57, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(57));
    
    \RDATA_IM_xhdl4[4]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_4, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(4));
    
    \curr_state[0]\ : SLE
      port map(D => N_384_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \curr_state[0]_net_1\);
    
    \RDATA_IM_xhdl4[1]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_1, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(1));
    
    \RDATA_IM_xhdl4[34]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_34, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(34));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \RDATA_IM_xhdl4[55]\ : SLE
      port map(D => i22_mux_2_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(55));
    
    \RDATA_IM_xhdl4[51]\ : SLE
      port map(D => N_8_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(51));
    
    \RDATA_IM_xhdl4[62]\ : SLE
      port map(D => i17_mux_0_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(62));
    
    \RDATA_IM_xhdl4[44]\ : SLE
      port map(D => N_3092_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(44));
    
    RLAST_IM_xhdl5_RNO : CFG3
      generic map(INIT => x"04")

      port map(A => \N_3167_i\, B => axi_state_0, C => N_3297, Y
         => COREAXI_0_AXImslave16_RLAST_m);
    
    \RDATA_IM_xhdl4[3]\ : SLE
      port map(D => N_3170_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(3));
    
    \RDATA_IM_xhdl4[20]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_20, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(20));
    
    \RDATA_IM_xhdl4[10]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_10, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(10));
    
    RVALID_IM_xhdl3 : SLE
      port map(D => rvalid_im_int_xhdl42_1, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RVALID_IM0\);
    
    \RDATA_IM_xhdl4[2]\ : SLE
      port map(D => N_39, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(2));
    
    RVALID_IM_r_RNIEGS81 : CFG3
      generic map(INIT => x"8F")

      port map(A => \RVALID_IM_r\, B => RREADY_MI0, C => 
        \curr_state[0]_net_1\, Y => \N_3167_i\);
    
    \RDATA_IM_xhdl4[56]\ : SLE
      port map(D => i22_mux_1_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(56));
    
    \RDATA_IM_xhdl4[52]\ : SLE
      port map(D => i22_mux_5_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(52));
    
    \RDATA_IM_xhdl4[33]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_33, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(33));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RDATA_IM_xhdl4[43]\ : SLE
      port map(D => \COREAXI_0_AXImslave16_RDATA_m[43]\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(43));
    
    \RDATA_IM_xhdl4[60]\ : SLE
      port map(D => i22_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(60));
    
    \RDATA_IM_xhdl4[24]\ : SLE
      port map(D => N_79_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(24));
    
    \RDATA_IM_xhdl4[14]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_14, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(14));
    
    \curr_state[5]\ : SLE
      port map(D => N_391_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \curr_state[5]_net_1\);
    
    \RDATA_IM_xhdl4[38]\ : SLE
      port map(D => N_3098_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(38));
    
    \RDATA_IM_xhdl4[48]\ : SLE
      port map(D => i17_mux_2_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(48));
    
    \RDATA_IM_xhdl4[39]\ : SLE
      port map(D => N_3096_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(39));
    
    \RDATA_IM_xhdl4[37]\ : SLE
      port map(D => N_3100_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(37));
    
    rvalid_im_int_xhdl42_1_0_a2_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \N_3167_i\, B => N_3163, Y => 
        rvalid_im_int_xhdl42_1);
    
    \RDATA_IM_xhdl4[49]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_49, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(49));
    
    \RDATA_IM_xhdl4[47]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_47, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(47));
    
    \RDATA_IM_xhdl4[50]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_50, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(50));
    
    \RDATA_IM_xhdl4[35]\ : SLE
      port map(D => N_3169_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(35));
    
    \RDATA_IM_xhdl4[31]\ : SLE
      port map(D => N_67_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(31));
    
    \RDATA_IM_xhdl4[23]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_23, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(23));
    
    \RDATA_IM_xhdl4[13]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_13, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(13));
    
    \RDATA_IM_xhdl4[0]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_0, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(0));
    
    \RDATA_IM_xhdl4[45]\ : SLE
      port map(D => N_3064_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(45));
    
    \RDATA_IM_xhdl4[41]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_41, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(41));
    
    \curr_state_RNO[0]\ : CFG4
      generic map(INIT => x"8ACF")

      port map(A => \curr_state[5]_net_1\, B => 
        \curr_state[0]_net_1\, C => N_3163, D => \N_3167_i\, Y
         => N_384_i);
    
    \RDATA_IM_xhdl4[28]\ : SLE
      port map(D => N_75_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(28));
    
    \RDATA_IM_xhdl4[18]\ : SLE
      port map(D => N_70_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(18));
    
    \RDATA_IM_xhdl4[54]\ : SLE
      port map(D => i22_mux_3_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(54));
    
    \RDATA_IM_xhdl4[6]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_6, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(6));
    
    \RDATA_IM_xhdl4[29]\ : SLE
      port map(D => N_69_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(29));
    
    \RDATA_IM_xhdl4[19]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_19, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(19));
    
    \RDATA_IM_xhdl4[7]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_7, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(7));
    
    \RDATA_IM_xhdl4[27]\ : SLE
      port map(D => N_76_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(27));
    
    \RDATA_IM_xhdl4[17]\ : SLE
      port map(D => N_71_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(17));
    
    \RDATA_IM_xhdl4[63]\ : SLE
      port map(D => i17_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(63));
    
    \RDATA_IM_xhdl4[36]\ : SLE
      port map(D => N_3102_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(36));
    
    \RDATA_IM_xhdl4[32]\ : SLE
      port map(D => N_3066_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(32));
    
    \RDATA_IM_xhdl4[9]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_9, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(9));
    
    \RDATA_IM_xhdl4[46]\ : SLE
      port map(D => \COREAXI_0_AXImslave16_RDATA_m[46]\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(46));
    
    \RDATA_IM_xhdl4[42]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_42, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(42));
    
    \RDATA_IM_xhdl4_RNO[46]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => COREAXI_0_AXImslave16_RDATA_3, B => 
        RDATA_reg_3, C => \N_3167_i\, D => N_74, Y => 
        \COREAXI_0_AXImslave16_RDATA_m[46]\);
    
    \RDATA_IM_xhdl4[25]\ : SLE
      port map(D => N_78_mux_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(25));
    
    \RDATA_IM_xhdl4[21]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_21, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(21));
    
    \RDATA_IM_xhdl4[15]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_15, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(15));
    
    \RDATA_IM_xhdl4[11]\ : SLE
      port map(D => COREAXI_0_AXImslave16_RDATA_m_11, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RDATA_IM0(11));
    
    \RDATA_IM_xhdl4_RNO[43]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => COREAXI_0_AXImslave16_RDATA_0, B => 
        RDATA_reg_0, C => \N_3167_i\, D => N_74, Y => 
        \COREAXI_0_AXImslave16_RDATA_m[43]\);
    
    RVALID_IM_r : SLE
      port map(D => \RVALID_IM0\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RVALID_IM_r\);
    
    RLAST_IM_xhdl5 : SLE
      port map(D => COREAXI_0_AXImslave16_RLAST_m, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => MSS_READY, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RLAST_IM0);
    
    \RDATA_IM_xhdl4[53]\ : SLE
      port map(D => i22_mux_4_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RDATA_IM0(53));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_rd_channel is

    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic;
          RDATA_reg_3                        : in    std_logic;
          RDATA_reg_0                        : in    std_logic;
          axi_state_0                        : in    std_logic;
          MSS_READY                          : in    std_logic;
          SDRCLK_c                           : in    std_logic;
          i22_mux_1_i                        : in    std_logic;
          i22_mux_0_i                        : in    std_logic;
          i22_mux_i                          : in    std_logic;
          i17_mux_1_i                        : in    std_logic;
          i17_mux_0_i                        : in    std_logic;
          i17_mux_i                          : in    std_logic;
          N_3092_i                           : in    std_logic;
          N_3064_i                           : in    std_logic;
          i17_mux_2_i                        : in    std_logic;
          N_8_i                              : in    std_logic;
          i22_mux_5_i                        : in    std_logic;
          i22_mux_4_i                        : in    std_logic;
          i22_mux_3_i                        : in    std_logic;
          i22_mux_2_i                        : in    std_logic;
          N_77_mux_i                         : in    std_logic;
          N_76_mux_i                         : in    std_logic;
          N_75_mux_i                         : in    std_logic;
          N_69_mux_i                         : in    std_logic;
          N_68_mux_i                         : in    std_logic;
          N_67_mux_i                         : in    std_logic;
          N_3066_i                           : in    std_logic;
          N_3169_i                           : in    std_logic;
          N_3102_i                           : in    std_logic;
          N_3100_i                           : in    std_logic;
          N_3098_i                           : in    std_logic;
          N_3096_i                           : in    std_logic;
          N_3094_i                           : in    std_logic;
          N_72_mux_i                         : in    std_logic;
          N_71_mux_i                         : in    std_logic;
          N_70_mux_i                         : in    std_logic;
          N_80_mux_i                         : in    std_logic;
          N_79_mux_i                         : in    std_logic;
          N_78_mux_i                         : in    std_logic;
          N_39                               : in    std_logic;
          N_3170_i                           : in    std_logic;
          RLAST_IM0                          : out   std_logic;
          RVALID_IM0                         : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic;
          N_23                               : out   std_logic;
          N_3167_i                           : out   std_logic;
          N_74                               : in    std_logic;
          N_389                              : in    std_logic;
          RREADY_MI0                         : in    std_logic;
          N_3297                             : in    std_logic
        );

end axi_rd_channel;

architecture DEF_ARCH of axi_rd_channel is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component axi_rdmatrix_16Sto1M
    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          axi_state_0                        : in    std_logic := 'U';
          RDATA_reg_3                        : in    std_logic := 'U';
          RDATA_reg_0                        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic := 'U';
          N_3297                             : in    std_logic := 'U';
          RREADY_MI0                         : in    std_logic := 'U';
          N_389                              : in    std_logic := 'U';
          N_74                               : in    std_logic := 'U';
          N_3167_i                           : out   std_logic;
          N_23                               : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic := 'U';
          RVALID_IM0                         : out   std_logic;
          RLAST_IM0                          : out   std_logic;
          N_3170_i                           : in    std_logic := 'U';
          N_39                               : in    std_logic := 'U';
          N_78_mux_i                         : in    std_logic := 'U';
          N_79_mux_i                         : in    std_logic := 'U';
          N_80_mux_i                         : in    std_logic := 'U';
          N_70_mux_i                         : in    std_logic := 'U';
          N_71_mux_i                         : in    std_logic := 'U';
          N_72_mux_i                         : in    std_logic := 'U';
          N_3094_i                           : in    std_logic := 'U';
          N_3096_i                           : in    std_logic := 'U';
          N_3098_i                           : in    std_logic := 'U';
          N_3100_i                           : in    std_logic := 'U';
          N_3102_i                           : in    std_logic := 'U';
          N_3169_i                           : in    std_logic := 'U';
          N_3066_i                           : in    std_logic := 'U';
          N_67_mux_i                         : in    std_logic := 'U';
          N_68_mux_i                         : in    std_logic := 'U';
          N_69_mux_i                         : in    std_logic := 'U';
          N_75_mux_i                         : in    std_logic := 'U';
          N_76_mux_i                         : in    std_logic := 'U';
          N_77_mux_i                         : in    std_logic := 'U';
          i22_mux_2_i                        : in    std_logic := 'U';
          i22_mux_3_i                        : in    std_logic := 'U';
          i22_mux_4_i                        : in    std_logic := 'U';
          i22_mux_5_i                        : in    std_logic := 'U';
          N_8_i                              : in    std_logic := 'U';
          i17_mux_2_i                        : in    std_logic := 'U';
          N_3064_i                           : in    std_logic := 'U';
          N_3092_i                           : in    std_logic := 'U';
          i17_mux_i                          : in    std_logic := 'U';
          i17_mux_0_i                        : in    std_logic := 'U';
          i17_mux_1_i                        : in    std_logic := 'U';
          i22_mux_i                          : in    std_logic := 'U';
          i22_mux_0_i                        : in    std_logic := 'U';
          i22_mux_1_i                        : in    std_logic := 'U';
          SDRCLK_c                           : in    std_logic := 'U';
          MSS_READY                          : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : axi_rdmatrix_16Sto1M
	Use entity work.axi_rdmatrix_16Sto1M(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    inst_rdmatrix_16Sto1M : axi_rdmatrix_16Sto1M
      port map(RDATA_IM0(63) => RDATA_IM0(63), RDATA_IM0(62) => 
        RDATA_IM0(62), RDATA_IM0(61) => RDATA_IM0(61), 
        RDATA_IM0(60) => RDATA_IM0(60), RDATA_IM0(59) => 
        RDATA_IM0(59), RDATA_IM0(58) => RDATA_IM0(58), 
        RDATA_IM0(57) => RDATA_IM0(57), RDATA_IM0(56) => 
        RDATA_IM0(56), RDATA_IM0(55) => RDATA_IM0(55), 
        RDATA_IM0(54) => RDATA_IM0(54), RDATA_IM0(53) => 
        RDATA_IM0(53), RDATA_IM0(52) => RDATA_IM0(52), 
        RDATA_IM0(51) => RDATA_IM0(51), RDATA_IM0(50) => 
        RDATA_IM0(50), RDATA_IM0(49) => RDATA_IM0(49), 
        RDATA_IM0(48) => RDATA_IM0(48), RDATA_IM0(47) => 
        RDATA_IM0(47), RDATA_IM0(46) => RDATA_IM0(46), 
        RDATA_IM0(45) => RDATA_IM0(45), RDATA_IM0(44) => 
        RDATA_IM0(44), RDATA_IM0(43) => RDATA_IM0(43), 
        RDATA_IM0(42) => RDATA_IM0(42), RDATA_IM0(41) => 
        RDATA_IM0(41), RDATA_IM0(40) => RDATA_IM0(40), 
        RDATA_IM0(39) => RDATA_IM0(39), RDATA_IM0(38) => 
        RDATA_IM0(38), RDATA_IM0(37) => RDATA_IM0(37), 
        RDATA_IM0(36) => RDATA_IM0(36), RDATA_IM0(35) => 
        RDATA_IM0(35), RDATA_IM0(34) => RDATA_IM0(34), 
        RDATA_IM0(33) => RDATA_IM0(33), RDATA_IM0(32) => 
        RDATA_IM0(32), RDATA_IM0(31) => RDATA_IM0(31), 
        RDATA_IM0(30) => RDATA_IM0(30), RDATA_IM0(29) => 
        RDATA_IM0(29), RDATA_IM0(28) => RDATA_IM0(28), 
        RDATA_IM0(27) => RDATA_IM0(27), RDATA_IM0(26) => 
        RDATA_IM0(26), RDATA_IM0(25) => RDATA_IM0(25), 
        RDATA_IM0(24) => RDATA_IM0(24), RDATA_IM0(23) => 
        RDATA_IM0(23), RDATA_IM0(22) => RDATA_IM0(22), 
        RDATA_IM0(21) => RDATA_IM0(21), RDATA_IM0(20) => 
        RDATA_IM0(20), RDATA_IM0(19) => RDATA_IM0(19), 
        RDATA_IM0(18) => RDATA_IM0(18), RDATA_IM0(17) => 
        RDATA_IM0(17), RDATA_IM0(16) => RDATA_IM0(16), 
        RDATA_IM0(15) => RDATA_IM0(15), RDATA_IM0(14) => 
        RDATA_IM0(14), RDATA_IM0(13) => RDATA_IM0(13), 
        RDATA_IM0(12) => RDATA_IM0(12), RDATA_IM0(11) => 
        RDATA_IM0(11), RDATA_IM0(10) => RDATA_IM0(10), 
        RDATA_IM0(9) => RDATA_IM0(9), RDATA_IM0(8) => 
        RDATA_IM0(8), RDATA_IM0(7) => RDATA_IM0(7), RDATA_IM0(6)
         => RDATA_IM0(6), RDATA_IM0(5) => RDATA_IM0(5), 
        RDATA_IM0(4) => RDATA_IM0(4), RDATA_IM0(3) => 
        RDATA_IM0(3), RDATA_IM0(2) => RDATA_IM0(2), RDATA_IM0(1)
         => RDATA_IM0(1), RDATA_IM0(0) => RDATA_IM0(0), 
        axi_state_0 => axi_state_0, RDATA_reg_3 => RDATA_reg_3, 
        RDATA_reg_0 => RDATA_reg_0, COREAXI_0_AXImslave16_RDATA_3
         => COREAXI_0_AXImslave16_RDATA_3, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        COREAXI_0_AXImslave16_RDATA_0, 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        COREAXI_0_AXImslave16_RDATA_m_57, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        COREAXI_0_AXImslave16_RDATA_m_58, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        COREAXI_0_AXImslave16_RDATA_m_41, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        COREAXI_0_AXImslave16_RDATA_m_42, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        COREAXI_0_AXImslave16_RDATA_m_47, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        COREAXI_0_AXImslave16_RDATA_m_49, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        COREAXI_0_AXImslave16_RDATA_m_50, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        COREAXI_0_AXImslave16_RDATA_m_33, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        COREAXI_0_AXImslave16_RDATA_m_34, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        COREAXI_0_AXImslave16_RDATA_m_11, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        COREAXI_0_AXImslave16_RDATA_m_12, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        COREAXI_0_AXImslave16_RDATA_m_13, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        COREAXI_0_AXImslave16_RDATA_m_14, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        COREAXI_0_AXImslave16_RDATA_m_15, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        COREAXI_0_AXImslave16_RDATA_m_19, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        COREAXI_0_AXImslave16_RDATA_m_20, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        COREAXI_0_AXImslave16_RDATA_m_21, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        COREAXI_0_AXImslave16_RDATA_m_23, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        COREAXI_0_AXImslave16_RDATA_m_0, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        COREAXI_0_AXImslave16_RDATA_m_1, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        COREAXI_0_AXImslave16_RDATA_m_4, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        COREAXI_0_AXImslave16_RDATA_m_5, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        COREAXI_0_AXImslave16_RDATA_m_6, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        COREAXI_0_AXImslave16_RDATA_m_7, 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        COREAXI_0_AXImslave16_RDATA_m_8, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        COREAXI_0_AXImslave16_RDATA_m_9, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        COREAXI_0_AXImslave16_RDATA_m_10, N_3297 => N_3297, 
        RREADY_MI0 => RREADY_MI0, N_389 => N_389, N_74 => N_74, 
        N_3167_i => N_3167_i, N_23 => N_23, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, RVALID_IM0 => 
        RVALID_IM0, RLAST_IM0 => RLAST_IM0, N_3170_i => N_3170_i, 
        N_39 => N_39, N_78_mux_i => N_78_mux_i, N_79_mux_i => 
        N_79_mux_i, N_80_mux_i => N_80_mux_i, N_70_mux_i => 
        N_70_mux_i, N_71_mux_i => N_71_mux_i, N_72_mux_i => 
        N_72_mux_i, N_3094_i => N_3094_i, N_3096_i => N_3096_i, 
        N_3098_i => N_3098_i, N_3100_i => N_3100_i, N_3102_i => 
        N_3102_i, N_3169_i => N_3169_i, N_3066_i => N_3066_i, 
        N_67_mux_i => N_67_mux_i, N_68_mux_i => N_68_mux_i, 
        N_69_mux_i => N_69_mux_i, N_75_mux_i => N_75_mux_i, 
        N_76_mux_i => N_76_mux_i, N_77_mux_i => N_77_mux_i, 
        i22_mux_2_i => i22_mux_2_i, i22_mux_3_i => i22_mux_3_i, 
        i22_mux_4_i => i22_mux_4_i, i22_mux_5_i => i22_mux_5_i, 
        N_8_i => N_8_i, i17_mux_2_i => i17_mux_2_i, N_3064_i => 
        N_3064_i, N_3092_i => N_3092_i, i17_mux_i => i17_mux_i, 
        i17_mux_0_i => i17_mux_0_i, i17_mux_1_i => i17_mux_1_i, 
        i22_mux_i => i22_mux_i, i22_mux_0_i => i22_mux_0_i, 
        i22_mux_1_i => i22_mux_1_i, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_wresp_channel is

    port( COREAXI_0_AXImslave16_BVALID : in    std_logic;
          SDRCLK_c                     : in    std_logic;
          MSS_READY                    : in    std_logic;
          BVALID_IM0                   : out   std_logic
        );

end axi_wresp_channel;

architecture DEF_ARCH of axi_wresp_channel is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    BVALID_IM_xhdl3 : SLE
      port map(D => COREAXI_0_AXImslave16_BVALID, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        BVALID_IM0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_matrix_m is

    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          axi_state_0                        : in    std_logic;
          RDATA_reg_3                        : in    std_logic;
          RDATA_reg_0                        : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic;
          BVALID_IM0                         : out   std_logic;
          COREAXI_0_AXImslave16_BVALID       : in    std_logic;
          N_3297                             : in    std_logic;
          RREADY_MI0                         : in    std_logic;
          N_389                              : in    std_logic;
          N_74                               : in    std_logic;
          N_3167_i                           : out   std_logic;
          N_23                               : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic;
          RVALID_IM0                         : out   std_logic;
          RLAST_IM0                          : out   std_logic;
          N_3170_i                           : in    std_logic;
          N_39                               : in    std_logic;
          N_78_mux_i                         : in    std_logic;
          N_79_mux_i                         : in    std_logic;
          N_80_mux_i                         : in    std_logic;
          N_70_mux_i                         : in    std_logic;
          N_71_mux_i                         : in    std_logic;
          N_72_mux_i                         : in    std_logic;
          N_3094_i                           : in    std_logic;
          N_3096_i                           : in    std_logic;
          N_3098_i                           : in    std_logic;
          N_3100_i                           : in    std_logic;
          N_3102_i                           : in    std_logic;
          N_3169_i                           : in    std_logic;
          N_3066_i                           : in    std_logic;
          N_67_mux_i                         : in    std_logic;
          N_68_mux_i                         : in    std_logic;
          N_69_mux_i                         : in    std_logic;
          N_75_mux_i                         : in    std_logic;
          N_76_mux_i                         : in    std_logic;
          N_77_mux_i                         : in    std_logic;
          i22_mux_2_i                        : in    std_logic;
          i22_mux_3_i                        : in    std_logic;
          i22_mux_4_i                        : in    std_logic;
          i22_mux_5_i                        : in    std_logic;
          N_8_i                              : in    std_logic;
          i17_mux_2_i                        : in    std_logic;
          N_3064_i                           : in    std_logic;
          N_3092_i                           : in    std_logic;
          i17_mux_i                          : in    std_logic;
          i17_mux_0_i                        : in    std_logic;
          i17_mux_1_i                        : in    std_logic;
          i22_mux_i                          : in    std_logic;
          i22_mux_0_i                        : in    std_logic;
          i22_mux_1_i                        : in    std_logic;
          SDRCLK_c                           : in    std_logic;
          MSS_READY                          : in    std_logic
        );

end axi_matrix_m;

architecture DEF_ARCH of axi_matrix_m is 

  component axi_rd_channel
    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic := 'U';
          RDATA_reg_3                        : in    std_logic := 'U';
          RDATA_reg_0                        : in    std_logic := 'U';
          axi_state_0                        : in    std_logic := 'U';
          MSS_READY                          : in    std_logic := 'U';
          SDRCLK_c                           : in    std_logic := 'U';
          i22_mux_1_i                        : in    std_logic := 'U';
          i22_mux_0_i                        : in    std_logic := 'U';
          i22_mux_i                          : in    std_logic := 'U';
          i17_mux_1_i                        : in    std_logic := 'U';
          i17_mux_0_i                        : in    std_logic := 'U';
          i17_mux_i                          : in    std_logic := 'U';
          N_3092_i                           : in    std_logic := 'U';
          N_3064_i                           : in    std_logic := 'U';
          i17_mux_2_i                        : in    std_logic := 'U';
          N_8_i                              : in    std_logic := 'U';
          i22_mux_5_i                        : in    std_logic := 'U';
          i22_mux_4_i                        : in    std_logic := 'U';
          i22_mux_3_i                        : in    std_logic := 'U';
          i22_mux_2_i                        : in    std_logic := 'U';
          N_77_mux_i                         : in    std_logic := 'U';
          N_76_mux_i                         : in    std_logic := 'U';
          N_75_mux_i                         : in    std_logic := 'U';
          N_69_mux_i                         : in    std_logic := 'U';
          N_68_mux_i                         : in    std_logic := 'U';
          N_67_mux_i                         : in    std_logic := 'U';
          N_3066_i                           : in    std_logic := 'U';
          N_3169_i                           : in    std_logic := 'U';
          N_3102_i                           : in    std_logic := 'U';
          N_3100_i                           : in    std_logic := 'U';
          N_3098_i                           : in    std_logic := 'U';
          N_3096_i                           : in    std_logic := 'U';
          N_3094_i                           : in    std_logic := 'U';
          N_72_mux_i                         : in    std_logic := 'U';
          N_71_mux_i                         : in    std_logic := 'U';
          N_70_mux_i                         : in    std_logic := 'U';
          N_80_mux_i                         : in    std_logic := 'U';
          N_79_mux_i                         : in    std_logic := 'U';
          N_78_mux_i                         : in    std_logic := 'U';
          N_39                               : in    std_logic := 'U';
          N_3170_i                           : in    std_logic := 'U';
          RLAST_IM0                          : out   std_logic;
          RVALID_IM0                         : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic := 'U';
          N_23                               : out   std_logic;
          N_3167_i                           : out   std_logic;
          N_74                               : in    std_logic := 'U';
          N_389                              : in    std_logic := 'U';
          RREADY_MI0                         : in    std_logic := 'U';
          N_3297                             : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component axi_wresp_channel
    port( COREAXI_0_AXImslave16_BVALID : in    std_logic := 'U';
          SDRCLK_c                     : in    std_logic := 'U';
          MSS_READY                    : in    std_logic := 'U';
          BVALID_IM0                   : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : axi_rd_channel
	Use entity work.axi_rd_channel(DEF_ARCH);
    for all : axi_wresp_channel
	Use entity work.axi_wresp_channel(DEF_ARCH);
begin 


    inst_rd_channel : axi_rd_channel
      port map(RDATA_IM0(63) => RDATA_IM0(63), RDATA_IM0(62) => 
        RDATA_IM0(62), RDATA_IM0(61) => RDATA_IM0(61), 
        RDATA_IM0(60) => RDATA_IM0(60), RDATA_IM0(59) => 
        RDATA_IM0(59), RDATA_IM0(58) => RDATA_IM0(58), 
        RDATA_IM0(57) => RDATA_IM0(57), RDATA_IM0(56) => 
        RDATA_IM0(56), RDATA_IM0(55) => RDATA_IM0(55), 
        RDATA_IM0(54) => RDATA_IM0(54), RDATA_IM0(53) => 
        RDATA_IM0(53), RDATA_IM0(52) => RDATA_IM0(52), 
        RDATA_IM0(51) => RDATA_IM0(51), RDATA_IM0(50) => 
        RDATA_IM0(50), RDATA_IM0(49) => RDATA_IM0(49), 
        RDATA_IM0(48) => RDATA_IM0(48), RDATA_IM0(47) => 
        RDATA_IM0(47), RDATA_IM0(46) => RDATA_IM0(46), 
        RDATA_IM0(45) => RDATA_IM0(45), RDATA_IM0(44) => 
        RDATA_IM0(44), RDATA_IM0(43) => RDATA_IM0(43), 
        RDATA_IM0(42) => RDATA_IM0(42), RDATA_IM0(41) => 
        RDATA_IM0(41), RDATA_IM0(40) => RDATA_IM0(40), 
        RDATA_IM0(39) => RDATA_IM0(39), RDATA_IM0(38) => 
        RDATA_IM0(38), RDATA_IM0(37) => RDATA_IM0(37), 
        RDATA_IM0(36) => RDATA_IM0(36), RDATA_IM0(35) => 
        RDATA_IM0(35), RDATA_IM0(34) => RDATA_IM0(34), 
        RDATA_IM0(33) => RDATA_IM0(33), RDATA_IM0(32) => 
        RDATA_IM0(32), RDATA_IM0(31) => RDATA_IM0(31), 
        RDATA_IM0(30) => RDATA_IM0(30), RDATA_IM0(29) => 
        RDATA_IM0(29), RDATA_IM0(28) => RDATA_IM0(28), 
        RDATA_IM0(27) => RDATA_IM0(27), RDATA_IM0(26) => 
        RDATA_IM0(26), RDATA_IM0(25) => RDATA_IM0(25), 
        RDATA_IM0(24) => RDATA_IM0(24), RDATA_IM0(23) => 
        RDATA_IM0(23), RDATA_IM0(22) => RDATA_IM0(22), 
        RDATA_IM0(21) => RDATA_IM0(21), RDATA_IM0(20) => 
        RDATA_IM0(20), RDATA_IM0(19) => RDATA_IM0(19), 
        RDATA_IM0(18) => RDATA_IM0(18), RDATA_IM0(17) => 
        RDATA_IM0(17), RDATA_IM0(16) => RDATA_IM0(16), 
        RDATA_IM0(15) => RDATA_IM0(15), RDATA_IM0(14) => 
        RDATA_IM0(14), RDATA_IM0(13) => RDATA_IM0(13), 
        RDATA_IM0(12) => RDATA_IM0(12), RDATA_IM0(11) => 
        RDATA_IM0(11), RDATA_IM0(10) => RDATA_IM0(10), 
        RDATA_IM0(9) => RDATA_IM0(9), RDATA_IM0(8) => 
        RDATA_IM0(8), RDATA_IM0(7) => RDATA_IM0(7), RDATA_IM0(6)
         => RDATA_IM0(6), RDATA_IM0(5) => RDATA_IM0(5), 
        RDATA_IM0(4) => RDATA_IM0(4), RDATA_IM0(3) => 
        RDATA_IM0(3), RDATA_IM0(2) => RDATA_IM0(2), RDATA_IM0(1)
         => RDATA_IM0(1), RDATA_IM0(0) => RDATA_IM0(0), 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        COREAXI_0_AXImslave16_RDATA_m_57, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        COREAXI_0_AXImslave16_RDATA_m_58, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        COREAXI_0_AXImslave16_RDATA_m_41, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        COREAXI_0_AXImslave16_RDATA_m_42, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        COREAXI_0_AXImslave16_RDATA_m_47, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        COREAXI_0_AXImslave16_RDATA_m_49, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        COREAXI_0_AXImslave16_RDATA_m_50, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        COREAXI_0_AXImslave16_RDATA_m_33, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        COREAXI_0_AXImslave16_RDATA_m_34, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        COREAXI_0_AXImslave16_RDATA_m_11, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        COREAXI_0_AXImslave16_RDATA_m_12, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        COREAXI_0_AXImslave16_RDATA_m_13, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        COREAXI_0_AXImslave16_RDATA_m_14, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        COREAXI_0_AXImslave16_RDATA_m_15, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        COREAXI_0_AXImslave16_RDATA_m_19, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        COREAXI_0_AXImslave16_RDATA_m_20, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        COREAXI_0_AXImslave16_RDATA_m_21, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        COREAXI_0_AXImslave16_RDATA_m_23, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        COREAXI_0_AXImslave16_RDATA_m_0, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        COREAXI_0_AXImslave16_RDATA_m_1, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        COREAXI_0_AXImslave16_RDATA_m_4, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        COREAXI_0_AXImslave16_RDATA_m_5, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        COREAXI_0_AXImslave16_RDATA_m_6, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        COREAXI_0_AXImslave16_RDATA_m_7, 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        COREAXI_0_AXImslave16_RDATA_m_8, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        COREAXI_0_AXImslave16_RDATA_m_9, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        COREAXI_0_AXImslave16_RDATA_m_10, 
        COREAXI_0_AXImslave16_RDATA_3 => 
        COREAXI_0_AXImslave16_RDATA_3, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        COREAXI_0_AXImslave16_RDATA_0, RDATA_reg_3 => RDATA_reg_3, 
        RDATA_reg_0 => RDATA_reg_0, axi_state_0 => axi_state_0, 
        MSS_READY => MSS_READY, SDRCLK_c => SDRCLK_c, i22_mux_1_i
         => i22_mux_1_i, i22_mux_0_i => i22_mux_0_i, i22_mux_i
         => i22_mux_i, i17_mux_1_i => i17_mux_1_i, i17_mux_0_i
         => i17_mux_0_i, i17_mux_i => i17_mux_i, N_3092_i => 
        N_3092_i, N_3064_i => N_3064_i, i17_mux_2_i => 
        i17_mux_2_i, N_8_i => N_8_i, i22_mux_5_i => i22_mux_5_i, 
        i22_mux_4_i => i22_mux_4_i, i22_mux_3_i => i22_mux_3_i, 
        i22_mux_2_i => i22_mux_2_i, N_77_mux_i => N_77_mux_i, 
        N_76_mux_i => N_76_mux_i, N_75_mux_i => N_75_mux_i, 
        N_69_mux_i => N_69_mux_i, N_68_mux_i => N_68_mux_i, 
        N_67_mux_i => N_67_mux_i, N_3066_i => N_3066_i, N_3169_i
         => N_3169_i, N_3102_i => N_3102_i, N_3100_i => N_3100_i, 
        N_3098_i => N_3098_i, N_3096_i => N_3096_i, N_3094_i => 
        N_3094_i, N_72_mux_i => N_72_mux_i, N_71_mux_i => 
        N_71_mux_i, N_70_mux_i => N_70_mux_i, N_80_mux_i => 
        N_80_mux_i, N_79_mux_i => N_79_mux_i, N_78_mux_i => 
        N_78_mux_i, N_39 => N_39, N_3170_i => N_3170_i, RLAST_IM0
         => RLAST_IM0, RVALID_IM0 => RVALID_IM0, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, N_23 => N_23, 
        N_3167_i => N_3167_i, N_74 => N_74, N_389 => N_389, 
        RREADY_MI0 => RREADY_MI0, N_3297 => N_3297);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    inst_wresp_channel : axi_wresp_channel
      port map(COREAXI_0_AXImslave16_BVALID => 
        COREAXI_0_AXImslave16_BVALID, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY, BVALID_IM0 => BVALID_IM0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity axi_interconnect_ntom is

    port( AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1);
          AWADDR_IS16_gated                    : out   std_logic_vector(23 downto 1);
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          WDATA_MI0                            : in    std_logic_vector(63 downto 0);
          WSTRB_MI0                            : in    std_logic_vector(7 downto 0);
          WDATA_IS16_gated                     : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated                     : out   std_logic_vector(7 downto 0);
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1);
          ARADDR_IS16_gated                    : out   std_logic_vector(23 downto 1);
          ARSIZE_MI0                           : in    std_logic_vector(1 downto 0);
          RDATA_IM0                            : out   std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          AWLOCK_MI0_i_0                       : in    std_logic;
          ARBURST_IS16_gated_0                 : out   std_logic;
          ARBURST_MI0_0                        : in    std_logic;
          ARLOCK_MI0_i_0                       : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_8      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_3        : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_0        : in    std_logic;
          RDATA_reg_3                          : in    std_logic;
          RDATA_reg_0                          : in    std_logic;
          axi_state_0                          : in    std_logic;
          AWREADY_IM0                          : out   std_logic;
          N_75_i                               : in    std_logic;
          AWVALID_MI0                          : in    std_logic;
          AWREADY_SI16                         : in    std_logic;
          m0_wr_end                            : in    std_logic;
          WREADY_SI16                          : in    std_logic;
          WVALID_MI0                           : in    std_logic;
          WREADY_IM0                           : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic;
          ARVALID_MI0                          : in    std_logic;
          m0_rd_end                            : in    std_logic;
          i22_mux_1_i                          : in    std_logic;
          i22_mux_0_i                          : in    std_logic;
          i22_mux_i                            : in    std_logic;
          i17_mux_1_i                          : in    std_logic;
          i17_mux_0_i                          : in    std_logic;
          i17_mux_i                            : in    std_logic;
          N_3092_i                             : in    std_logic;
          N_3064_i                             : in    std_logic;
          i17_mux_2_i                          : in    std_logic;
          N_8_i                                : in    std_logic;
          i22_mux_5_i                          : in    std_logic;
          i22_mux_4_i                          : in    std_logic;
          i22_mux_3_i                          : in    std_logic;
          i22_mux_2_i                          : in    std_logic;
          N_77_mux_i                           : in    std_logic;
          N_76_mux_i                           : in    std_logic;
          N_75_mux_i                           : in    std_logic;
          N_69_mux_i                           : in    std_logic;
          N_68_mux_i                           : in    std_logic;
          N_67_mux_i                           : in    std_logic;
          N_3066_i                             : in    std_logic;
          N_3169_i                             : in    std_logic;
          N_3102_i                             : in    std_logic;
          N_3100_i                             : in    std_logic;
          N_3098_i                             : in    std_logic;
          N_3096_i                             : in    std_logic;
          N_3094_i                             : in    std_logic;
          N_72_mux_i                           : in    std_logic;
          N_71_mux_i                           : in    std_logic;
          N_70_mux_i                           : in    std_logic;
          N_80_mux_i                           : in    std_logic;
          N_79_mux_i                           : in    std_logic;
          N_78_mux_i                           : in    std_logic;
          N_39                                 : in    std_logic;
          N_3170_i                             : in    std_logic;
          RLAST_IM0                            : out   std_logic;
          RVALID_IM0                           : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic;
          N_23                                 : out   std_logic;
          N_3167_i                             : out   std_logic;
          N_74                                 : in    std_logic;
          N_389                                : in    std_logic;
          RREADY_MI0                           : in    std_logic;
          N_3297                               : in    std_logic;
          COREAXI_0_AXImslave16_BVALID         : in    std_logic;
          BVALID_IM0                           : out   std_logic;
          ARVALID_IS16                         : out   std_logic;
          AWVALID_IS16                         : out   std_logic;
          WVALID_IS16                          : out   std_logic;
          SDRCLK_c                             : in    std_logic;
          MSS_READY                            : in    std_logic
        );

end axi_interconnect_ntom;

architecture DEF_ARCH of axi_interconnect_ntom is 

  component axi_matrix_s
    port( ARSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          ARADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          WSTRB_IS16_gated                     : out   std_logic_vector(7 downto 0);
          WDATA_IS16_gated                     : out   std_logic_vector(63 downto 0);
          WSTRB_MI0                            : in    std_logic_vector(7 downto 0) := (others => 'U');
          WDATA_MI0                            : in    std_logic_vector(63 downto 0) := (others => 'U');
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          AWADDR_IS16_gated                    : out   std_logic_vector(27 downto 1);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARLOCK_MI0_i_0                       : in    std_logic := 'U';
          ARBURST_MI0_0                        : in    std_logic := 'U';
          ARBURST_IS16_gated_0                 : out   std_logic;
          AWLOCK_MI0_i_0                       : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          m0_rd_end                            : in    std_logic := 'U';
          ARVALID_MI0                          : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          ARVALID_IS16_gated                   : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          WREADY_IM0                           : out   std_logic;
          WVALID_IS16_gated                    : out   std_logic;
          WVALID_MI0                           : in    std_logic := 'U';
          WREADY_SI16                          : in    std_logic := 'U';
          m0_wr_end                            : in    std_logic := 'U';
          AWREADY_SI16                         : in    std_logic := 'U';
          AWVALID_MI0                          : in    std_logic := 'U';
          N_75_i                               : in    std_logic := 'U';
          AWVALID_IS16_gated                   : out   std_logic;
          AWREADY_IM0                          : out   std_logic;
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component axi_matrix_m
    port( RDATA_IM0                          : out   std_logic_vector(63 downto 0);
          axi_state_0                        : in    std_logic := 'U';
          RDATA_reg_3                        : in    std_logic := 'U';
          RDATA_reg_0                        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_3      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_0      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_57   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_58   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_41   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_42   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_47   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_49   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_50   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_33   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_34   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_11   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_12   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_13   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_14   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_15   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_19   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_20   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_21   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_23   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_0    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_1    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_4    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_5    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_6    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_7    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_8    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_9    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_10   : in    std_logic := 'U';
          BVALID_IM0                         : out   std_logic;
          COREAXI_0_AXImslave16_BVALID       : in    std_logic := 'U';
          N_3297                             : in    std_logic := 'U';
          RREADY_MI0                         : in    std_logic := 'U';
          N_389                              : in    std_logic := 'U';
          N_74                               : in    std_logic := 'U';
          N_3167_i                           : out   std_logic;
          N_23                               : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RREADY : in    std_logic := 'U';
          RVALID_IM0                         : out   std_logic;
          RLAST_IM0                          : out   std_logic;
          N_3170_i                           : in    std_logic := 'U';
          N_39                               : in    std_logic := 'U';
          N_78_mux_i                         : in    std_logic := 'U';
          N_79_mux_i                         : in    std_logic := 'U';
          N_80_mux_i                         : in    std_logic := 'U';
          N_70_mux_i                         : in    std_logic := 'U';
          N_71_mux_i                         : in    std_logic := 'U';
          N_72_mux_i                         : in    std_logic := 'U';
          N_3094_i                           : in    std_logic := 'U';
          N_3096_i                           : in    std_logic := 'U';
          N_3098_i                           : in    std_logic := 'U';
          N_3100_i                           : in    std_logic := 'U';
          N_3102_i                           : in    std_logic := 'U';
          N_3169_i                           : in    std_logic := 'U';
          N_3066_i                           : in    std_logic := 'U';
          N_67_mux_i                         : in    std_logic := 'U';
          N_68_mux_i                         : in    std_logic := 'U';
          N_69_mux_i                         : in    std_logic := 'U';
          N_75_mux_i                         : in    std_logic := 'U';
          N_76_mux_i                         : in    std_logic := 'U';
          N_77_mux_i                         : in    std_logic := 'U';
          i22_mux_2_i                        : in    std_logic := 'U';
          i22_mux_3_i                        : in    std_logic := 'U';
          i22_mux_4_i                        : in    std_logic := 'U';
          i22_mux_5_i                        : in    std_logic := 'U';
          N_8_i                              : in    std_logic := 'U';
          i17_mux_2_i                        : in    std_logic := 'U';
          N_3064_i                           : in    std_logic := 'U';
          N_3092_i                           : in    std_logic := 'U';
          i17_mux_i                          : in    std_logic := 'U';
          i17_mux_0_i                        : in    std_logic := 'U';
          i17_mux_1_i                        : in    std_logic := 'U';
          i22_mux_i                          : in    std_logic := 'U';
          i22_mux_0_i                        : in    std_logic := 'U';
          i22_mux_1_i                        : in    std_logic := 'U';
          SDRCLK_c                           : in    std_logic := 'U';
          MSS_READY                          : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \ARADDR_IS16_gated_r[26]_net_1\, VCC_net_1, 
        \ARADDR_IS16_gated[26]\, GND_net_1, 
        \ARADDR_IS16_gated_r[27]_net_1\, \ARADDR_IS16_gated[27]\, 
        \AWADDR_IS16_gated_r[26]_net_1\, \AWADDR_IS16_gated[26]\, 
        \AWADDR_IS16_gated_r[27]_net_1\, \AWADDR_IS16_gated[27]\, 
        \AWVALID_IS16_gated_r\, AWVALID_IS16_gated, 
        \WVALID_IS16_gated_r\, WVALID_IS16_gated, 
        \ARVALID_IS16_gated_r\, ARVALID_IS16_gated : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

    for all : axi_matrix_s
	Use entity work.axi_matrix_s(DEF_ARCH);
    for all : axi_matrix_m
	Use entity work.axi_matrix_m(DEF_ARCH);
begin 


    \L27.inst_matrix_S16\ : axi_matrix_s
      port map(ARSIZE_MI0(1) => ARSIZE_MI0(1), ARSIZE_MI0(0) => 
        ARSIZE_MI0(0), ARADDR_IS16_gated(27) => 
        \ARADDR_IS16_gated[27]\, ARADDR_IS16_gated(26) => 
        \ARADDR_IS16_gated[26]\, ARADDR_IS16_gated(25) => nc8, 
        ARADDR_IS16_gated(24) => nc7, ARADDR_IS16_gated(23) => 
        ARADDR_IS16_gated(23), ARADDR_IS16_gated(22) => 
        ARADDR_IS16_gated(22), ARADDR_IS16_gated(21) => 
        ARADDR_IS16_gated(21), ARADDR_IS16_gated(20) => 
        ARADDR_IS16_gated(20), ARADDR_IS16_gated(19) => 
        ARADDR_IS16_gated(19), ARADDR_IS16_gated(18) => 
        ARADDR_IS16_gated(18), ARADDR_IS16_gated(17) => 
        ARADDR_IS16_gated(17), ARADDR_IS16_gated(16) => 
        ARADDR_IS16_gated(16), ARADDR_IS16_gated(15) => 
        ARADDR_IS16_gated(15), ARADDR_IS16_gated(14) => 
        ARADDR_IS16_gated(14), ARADDR_IS16_gated(13) => 
        ARADDR_IS16_gated(13), ARADDR_IS16_gated(12) => 
        ARADDR_IS16_gated(12), ARADDR_IS16_gated(11) => 
        ARADDR_IS16_gated(11), ARADDR_IS16_gated(10) => 
        ARADDR_IS16_gated(10), ARADDR_IS16_gated(9) => 
        ARADDR_IS16_gated(9), ARADDR_IS16_gated(8) => 
        ARADDR_IS16_gated(8), ARADDR_IS16_gated(7) => 
        ARADDR_IS16_gated(7), ARADDR_IS16_gated(6) => 
        ARADDR_IS16_gated(6), ARADDR_IS16_gated(5) => 
        ARADDR_IS16_gated(5), ARADDR_IS16_gated(4) => 
        ARADDR_IS16_gated(4), ARADDR_IS16_gated(3) => 
        ARADDR_IS16_gated(3), ARADDR_IS16_gated(2) => 
        ARADDR_IS16_gated(2), ARADDR_IS16_gated(1) => 
        ARADDR_IS16_gated(1), ARADDR_MI0(27) => ARADDR_MI0(27), 
        ARADDR_MI0(26) => ARADDR_MI0(26), ARADDR_MI0(25) => nc6, 
        ARADDR_MI0(24) => nc2, ARADDR_MI0(23) => ARADDR_MI0(23), 
        ARADDR_MI0(22) => ARADDR_MI0(22), ARADDR_MI0(21) => 
        ARADDR_MI0(21), ARADDR_MI0(20) => ARADDR_MI0(20), 
        ARADDR_MI0(19) => ARADDR_MI0(19), ARADDR_MI0(18) => 
        ARADDR_MI0(18), ARADDR_MI0(17) => ARADDR_MI0(17), 
        ARADDR_MI0(16) => ARADDR_MI0(16), ARADDR_MI0(15) => 
        ARADDR_MI0(15), ARADDR_MI0(14) => ARADDR_MI0(14), 
        ARADDR_MI0(13) => ARADDR_MI0(13), ARADDR_MI0(12) => 
        ARADDR_MI0(12), ARADDR_MI0(11) => ARADDR_MI0(11), 
        ARADDR_MI0(10) => ARADDR_MI0(10), ARADDR_MI0(9) => 
        ARADDR_MI0(9), ARADDR_MI0(8) => ARADDR_MI0(8), 
        ARADDR_MI0(7) => ARADDR_MI0(7), ARADDR_MI0(6) => 
        ARADDR_MI0(6), ARADDR_MI0(5) => ARADDR_MI0(5), 
        ARADDR_MI0(4) => ARADDR_MI0(4), ARADDR_MI0(3) => 
        ARADDR_MI0(3), ARADDR_MI0(2) => ARADDR_MI0(2), 
        ARADDR_MI0(1) => ARADDR_MI0(1), ARSIZE_IS16_gated(1) => 
        ARSIZE_IS16_gated(1), ARSIZE_IS16_gated(0) => 
        ARSIZE_IS16_gated(0), WSTRB_IS16_gated(7) => 
        WSTRB_IS16_gated(7), WSTRB_IS16_gated(6) => 
        WSTRB_IS16_gated(6), WSTRB_IS16_gated(5) => 
        WSTRB_IS16_gated(5), WSTRB_IS16_gated(4) => 
        WSTRB_IS16_gated(4), WSTRB_IS16_gated(3) => 
        WSTRB_IS16_gated(3), WSTRB_IS16_gated(2) => 
        WSTRB_IS16_gated(2), WSTRB_IS16_gated(1) => 
        WSTRB_IS16_gated(1), WSTRB_IS16_gated(0) => 
        WSTRB_IS16_gated(0), WDATA_IS16_gated(63) => 
        WDATA_IS16_gated(63), WDATA_IS16_gated(62) => 
        WDATA_IS16_gated(62), WDATA_IS16_gated(61) => 
        WDATA_IS16_gated(61), WDATA_IS16_gated(60) => 
        WDATA_IS16_gated(60), WDATA_IS16_gated(59) => 
        WDATA_IS16_gated(59), WDATA_IS16_gated(58) => 
        WDATA_IS16_gated(58), WDATA_IS16_gated(57) => 
        WDATA_IS16_gated(57), WDATA_IS16_gated(56) => 
        WDATA_IS16_gated(56), WDATA_IS16_gated(55) => 
        WDATA_IS16_gated(55), WDATA_IS16_gated(54) => 
        WDATA_IS16_gated(54), WDATA_IS16_gated(53) => 
        WDATA_IS16_gated(53), WDATA_IS16_gated(52) => 
        WDATA_IS16_gated(52), WDATA_IS16_gated(51) => 
        WDATA_IS16_gated(51), WDATA_IS16_gated(50) => 
        WDATA_IS16_gated(50), WDATA_IS16_gated(49) => 
        WDATA_IS16_gated(49), WDATA_IS16_gated(48) => 
        WDATA_IS16_gated(48), WDATA_IS16_gated(47) => 
        WDATA_IS16_gated(47), WDATA_IS16_gated(46) => 
        WDATA_IS16_gated(46), WDATA_IS16_gated(45) => 
        WDATA_IS16_gated(45), WDATA_IS16_gated(44) => 
        WDATA_IS16_gated(44), WDATA_IS16_gated(43) => 
        WDATA_IS16_gated(43), WDATA_IS16_gated(42) => 
        WDATA_IS16_gated(42), WDATA_IS16_gated(41) => 
        WDATA_IS16_gated(41), WDATA_IS16_gated(40) => 
        WDATA_IS16_gated(40), WDATA_IS16_gated(39) => 
        WDATA_IS16_gated(39), WDATA_IS16_gated(38) => 
        WDATA_IS16_gated(38), WDATA_IS16_gated(37) => 
        WDATA_IS16_gated(37), WDATA_IS16_gated(36) => 
        WDATA_IS16_gated(36), WDATA_IS16_gated(35) => 
        WDATA_IS16_gated(35), WDATA_IS16_gated(34) => 
        WDATA_IS16_gated(34), WDATA_IS16_gated(33) => 
        WDATA_IS16_gated(33), WDATA_IS16_gated(32) => 
        WDATA_IS16_gated(32), WDATA_IS16_gated(31) => 
        WDATA_IS16_gated(31), WDATA_IS16_gated(30) => 
        WDATA_IS16_gated(30), WDATA_IS16_gated(29) => 
        WDATA_IS16_gated(29), WDATA_IS16_gated(28) => 
        WDATA_IS16_gated(28), WDATA_IS16_gated(27) => 
        WDATA_IS16_gated(27), WDATA_IS16_gated(26) => 
        WDATA_IS16_gated(26), WDATA_IS16_gated(25) => 
        WDATA_IS16_gated(25), WDATA_IS16_gated(24) => 
        WDATA_IS16_gated(24), WDATA_IS16_gated(23) => 
        WDATA_IS16_gated(23), WDATA_IS16_gated(22) => 
        WDATA_IS16_gated(22), WDATA_IS16_gated(21) => 
        WDATA_IS16_gated(21), WDATA_IS16_gated(20) => 
        WDATA_IS16_gated(20), WDATA_IS16_gated(19) => 
        WDATA_IS16_gated(19), WDATA_IS16_gated(18) => 
        WDATA_IS16_gated(18), WDATA_IS16_gated(17) => 
        WDATA_IS16_gated(17), WDATA_IS16_gated(16) => 
        WDATA_IS16_gated(16), WDATA_IS16_gated(15) => 
        WDATA_IS16_gated(15), WDATA_IS16_gated(14) => 
        WDATA_IS16_gated(14), WDATA_IS16_gated(13) => 
        WDATA_IS16_gated(13), WDATA_IS16_gated(12) => 
        WDATA_IS16_gated(12), WDATA_IS16_gated(11) => 
        WDATA_IS16_gated(11), WDATA_IS16_gated(10) => 
        WDATA_IS16_gated(10), WDATA_IS16_gated(9) => 
        WDATA_IS16_gated(9), WDATA_IS16_gated(8) => 
        WDATA_IS16_gated(8), WDATA_IS16_gated(7) => 
        WDATA_IS16_gated(7), WDATA_IS16_gated(6) => 
        WDATA_IS16_gated(6), WDATA_IS16_gated(5) => 
        WDATA_IS16_gated(5), WDATA_IS16_gated(4) => 
        WDATA_IS16_gated(4), WDATA_IS16_gated(3) => 
        WDATA_IS16_gated(3), WDATA_IS16_gated(2) => 
        WDATA_IS16_gated(2), WDATA_IS16_gated(1) => 
        WDATA_IS16_gated(1), WDATA_IS16_gated(0) => 
        WDATA_IS16_gated(0), WSTRB_MI0(7) => WSTRB_MI0(7), 
        WSTRB_MI0(6) => WSTRB_MI0(6), WSTRB_MI0(5) => 
        WSTRB_MI0(5), WSTRB_MI0(4) => WSTRB_MI0(4), WSTRB_MI0(3)
         => WSTRB_MI0(3), WSTRB_MI0(2) => WSTRB_MI0(2), 
        WSTRB_MI0(1) => WSTRB_MI0(1), WSTRB_MI0(0) => 
        WSTRB_MI0(0), WDATA_MI0(63) => WDATA_MI0(63), 
        WDATA_MI0(62) => WDATA_MI0(62), WDATA_MI0(61) => 
        WDATA_MI0(61), WDATA_MI0(60) => WDATA_MI0(60), 
        WDATA_MI0(59) => WDATA_MI0(59), WDATA_MI0(58) => 
        WDATA_MI0(58), WDATA_MI0(57) => WDATA_MI0(57), 
        WDATA_MI0(56) => WDATA_MI0(56), WDATA_MI0(55) => 
        WDATA_MI0(55), WDATA_MI0(54) => WDATA_MI0(54), 
        WDATA_MI0(53) => WDATA_MI0(53), WDATA_MI0(52) => 
        WDATA_MI0(52), WDATA_MI0(51) => WDATA_MI0(51), 
        WDATA_MI0(50) => WDATA_MI0(50), WDATA_MI0(49) => 
        WDATA_MI0(49), WDATA_MI0(48) => WDATA_MI0(48), 
        WDATA_MI0(47) => WDATA_MI0(47), WDATA_MI0(46) => 
        WDATA_MI0(46), WDATA_MI0(45) => WDATA_MI0(45), 
        WDATA_MI0(44) => WDATA_MI0(44), WDATA_MI0(43) => 
        WDATA_MI0(43), WDATA_MI0(42) => WDATA_MI0(42), 
        WDATA_MI0(41) => WDATA_MI0(41), WDATA_MI0(40) => 
        WDATA_MI0(40), WDATA_MI0(39) => WDATA_MI0(39), 
        WDATA_MI0(38) => WDATA_MI0(38), WDATA_MI0(37) => 
        WDATA_MI0(37), WDATA_MI0(36) => WDATA_MI0(36), 
        WDATA_MI0(35) => WDATA_MI0(35), WDATA_MI0(34) => 
        WDATA_MI0(34), WDATA_MI0(33) => WDATA_MI0(33), 
        WDATA_MI0(32) => WDATA_MI0(32), WDATA_MI0(31) => 
        WDATA_MI0(31), WDATA_MI0(30) => WDATA_MI0(30), 
        WDATA_MI0(29) => WDATA_MI0(29), WDATA_MI0(28) => 
        WDATA_MI0(28), WDATA_MI0(27) => WDATA_MI0(27), 
        WDATA_MI0(26) => WDATA_MI0(26), WDATA_MI0(25) => 
        WDATA_MI0(25), WDATA_MI0(24) => WDATA_MI0(24), 
        WDATA_MI0(23) => WDATA_MI0(23), WDATA_MI0(22) => 
        WDATA_MI0(22), WDATA_MI0(21) => WDATA_MI0(21), 
        WDATA_MI0(20) => WDATA_MI0(20), WDATA_MI0(19) => 
        WDATA_MI0(19), WDATA_MI0(18) => WDATA_MI0(18), 
        WDATA_MI0(17) => WDATA_MI0(17), WDATA_MI0(16) => 
        WDATA_MI0(16), WDATA_MI0(15) => WDATA_MI0(15), 
        WDATA_MI0(14) => WDATA_MI0(14), WDATA_MI0(13) => 
        WDATA_MI0(13), WDATA_MI0(12) => WDATA_MI0(12), 
        WDATA_MI0(11) => WDATA_MI0(11), WDATA_MI0(10) => 
        WDATA_MI0(10), WDATA_MI0(9) => WDATA_MI0(9), WDATA_MI0(8)
         => WDATA_MI0(8), WDATA_MI0(7) => WDATA_MI0(7), 
        WDATA_MI0(6) => WDATA_MI0(6), WDATA_MI0(5) => 
        WDATA_MI0(5), WDATA_MI0(4) => WDATA_MI0(4), WDATA_MI0(3)
         => WDATA_MI0(3), WDATA_MI0(2) => WDATA_MI0(2), 
        WDATA_MI0(1) => WDATA_MI0(1), WDATA_MI0(0) => 
        WDATA_MI0(0), AWSIZE_MI0(1) => AWSIZE_MI0(1), 
        AWSIZE_MI0(0) => AWSIZE_MI0(0), AWADDR_IS16_gated(27) => 
        \AWADDR_IS16_gated[27]\, AWADDR_IS16_gated(26) => 
        \AWADDR_IS16_gated[26]\, AWADDR_IS16_gated(25) => nc5, 
        AWADDR_IS16_gated(24) => nc4, AWADDR_IS16_gated(23) => 
        AWADDR_IS16_gated(23), AWADDR_IS16_gated(22) => 
        AWADDR_IS16_gated(22), AWADDR_IS16_gated(21) => 
        AWADDR_IS16_gated(21), AWADDR_IS16_gated(20) => 
        AWADDR_IS16_gated(20), AWADDR_IS16_gated(19) => 
        AWADDR_IS16_gated(19), AWADDR_IS16_gated(18) => 
        AWADDR_IS16_gated(18), AWADDR_IS16_gated(17) => 
        AWADDR_IS16_gated(17), AWADDR_IS16_gated(16) => 
        AWADDR_IS16_gated(16), AWADDR_IS16_gated(15) => 
        AWADDR_IS16_gated(15), AWADDR_IS16_gated(14) => 
        AWADDR_IS16_gated(14), AWADDR_IS16_gated(13) => 
        AWADDR_IS16_gated(13), AWADDR_IS16_gated(12) => 
        AWADDR_IS16_gated(12), AWADDR_IS16_gated(11) => 
        AWADDR_IS16_gated(11), AWADDR_IS16_gated(10) => 
        AWADDR_IS16_gated(10), AWADDR_IS16_gated(9) => 
        AWADDR_IS16_gated(9), AWADDR_IS16_gated(8) => 
        AWADDR_IS16_gated(8), AWADDR_IS16_gated(7) => 
        AWADDR_IS16_gated(7), AWADDR_IS16_gated(6) => 
        AWADDR_IS16_gated(6), AWADDR_IS16_gated(5) => 
        AWADDR_IS16_gated(5), AWADDR_IS16_gated(4) => 
        AWADDR_IS16_gated(4), AWADDR_IS16_gated(3) => 
        AWADDR_IS16_gated(3), AWADDR_IS16_gated(2) => 
        AWADDR_IS16_gated(2), AWADDR_IS16_gated(1) => 
        AWADDR_IS16_gated(1), AWADDR_MI0(27) => AWADDR_MI0(27), 
        AWADDR_MI0(26) => AWADDR_MI0(26), AWADDR_MI0(25) => nc3, 
        AWADDR_MI0(24) => nc1, AWADDR_MI0(23) => AWADDR_MI0(23), 
        AWADDR_MI0(22) => AWADDR_MI0(22), AWADDR_MI0(21) => 
        AWADDR_MI0(21), AWADDR_MI0(20) => AWADDR_MI0(20), 
        AWADDR_MI0(19) => AWADDR_MI0(19), AWADDR_MI0(18) => 
        AWADDR_MI0(18), AWADDR_MI0(17) => AWADDR_MI0(17), 
        AWADDR_MI0(16) => AWADDR_MI0(16), AWADDR_MI0(15) => 
        AWADDR_MI0(15), AWADDR_MI0(14) => AWADDR_MI0(14), 
        AWADDR_MI0(13) => AWADDR_MI0(13), AWADDR_MI0(12) => 
        AWADDR_MI0(12), AWADDR_MI0(11) => AWADDR_MI0(11), 
        AWADDR_MI0(10) => AWADDR_MI0(10), AWADDR_MI0(9) => 
        AWADDR_MI0(9), AWADDR_MI0(8) => AWADDR_MI0(8), 
        AWADDR_MI0(7) => AWADDR_MI0(7), AWADDR_MI0(6) => 
        AWADDR_MI0(6), AWADDR_MI0(5) => AWADDR_MI0(5), 
        AWADDR_MI0(4) => AWADDR_MI0(4), AWADDR_MI0(3) => 
        AWADDR_MI0(3), AWADDR_MI0(2) => AWADDR_MI0(2), 
        AWADDR_MI0(1) => AWADDR_MI0(1), AWSIZE_IS16_gated(1) => 
        AWSIZE_IS16_gated(1), AWSIZE_IS16_gated(0) => 
        AWSIZE_IS16_gated(0), ARLOCK_MI0_i_0 => ARLOCK_MI0_i_0, 
        ARBURST_MI0_0 => ARBURST_MI0_0, ARBURST_IS16_gated_0 => 
        ARBURST_IS16_gated_0, AWLOCK_MI0_i_0 => AWLOCK_MI0_i_0, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, m0_rd_end => 
        m0_rd_end, ARVALID_MI0 => ARVALID_MI0, 
        COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, 
        COREAXI_0_AXImslave16_ARVALID => 
        COREAXI_0_AXImslave16_ARVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, ARVALID_IS16_gated
         => ARVALID_IS16_gated, ARREADY_IM0 => ARREADY_IM0, 
        WREADY_IM0 => WREADY_IM0, WVALID_IS16_gated => 
        WVALID_IS16_gated, WVALID_MI0 => WVALID_MI0, WREADY_SI16
         => WREADY_SI16, m0_wr_end => m0_wr_end, AWREADY_SI16 => 
        AWREADY_SI16, AWVALID_MI0 => AWVALID_MI0, N_75_i => 
        N_75_i, AWVALID_IS16_gated => AWVALID_IS16_gated, 
        AWREADY_IM0 => AWREADY_IM0, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY);
    
    ARVALID_IS16_gated_r : SLE
      port map(D => ARVALID_IS16_gated, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARVALID_IS16_gated_r\);
    
    \ARADDR_IS16_gated_r[26]\ : SLE
      port map(D => \ARADDR_IS16_gated[26]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS16_gated_r[26]_net_1\);
    
    \AWADDR_IS16_gated_r[26]\ : SLE
      port map(D => \AWADDR_IS16_gated[26]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWADDR_IS16_gated_r[26]_net_1\);
    
    inst_matrix_m0 : axi_matrix_m
      port map(RDATA_IM0(63) => RDATA_IM0(63), RDATA_IM0(62) => 
        RDATA_IM0(62), RDATA_IM0(61) => RDATA_IM0(61), 
        RDATA_IM0(60) => RDATA_IM0(60), RDATA_IM0(59) => 
        RDATA_IM0(59), RDATA_IM0(58) => RDATA_IM0(58), 
        RDATA_IM0(57) => RDATA_IM0(57), RDATA_IM0(56) => 
        RDATA_IM0(56), RDATA_IM0(55) => RDATA_IM0(55), 
        RDATA_IM0(54) => RDATA_IM0(54), RDATA_IM0(53) => 
        RDATA_IM0(53), RDATA_IM0(52) => RDATA_IM0(52), 
        RDATA_IM0(51) => RDATA_IM0(51), RDATA_IM0(50) => 
        RDATA_IM0(50), RDATA_IM0(49) => RDATA_IM0(49), 
        RDATA_IM0(48) => RDATA_IM0(48), RDATA_IM0(47) => 
        RDATA_IM0(47), RDATA_IM0(46) => RDATA_IM0(46), 
        RDATA_IM0(45) => RDATA_IM0(45), RDATA_IM0(44) => 
        RDATA_IM0(44), RDATA_IM0(43) => RDATA_IM0(43), 
        RDATA_IM0(42) => RDATA_IM0(42), RDATA_IM0(41) => 
        RDATA_IM0(41), RDATA_IM0(40) => RDATA_IM0(40), 
        RDATA_IM0(39) => RDATA_IM0(39), RDATA_IM0(38) => 
        RDATA_IM0(38), RDATA_IM0(37) => RDATA_IM0(37), 
        RDATA_IM0(36) => RDATA_IM0(36), RDATA_IM0(35) => 
        RDATA_IM0(35), RDATA_IM0(34) => RDATA_IM0(34), 
        RDATA_IM0(33) => RDATA_IM0(33), RDATA_IM0(32) => 
        RDATA_IM0(32), RDATA_IM0(31) => RDATA_IM0(31), 
        RDATA_IM0(30) => RDATA_IM0(30), RDATA_IM0(29) => 
        RDATA_IM0(29), RDATA_IM0(28) => RDATA_IM0(28), 
        RDATA_IM0(27) => RDATA_IM0(27), RDATA_IM0(26) => 
        RDATA_IM0(26), RDATA_IM0(25) => RDATA_IM0(25), 
        RDATA_IM0(24) => RDATA_IM0(24), RDATA_IM0(23) => 
        RDATA_IM0(23), RDATA_IM0(22) => RDATA_IM0(22), 
        RDATA_IM0(21) => RDATA_IM0(21), RDATA_IM0(20) => 
        RDATA_IM0(20), RDATA_IM0(19) => RDATA_IM0(19), 
        RDATA_IM0(18) => RDATA_IM0(18), RDATA_IM0(17) => 
        RDATA_IM0(17), RDATA_IM0(16) => RDATA_IM0(16), 
        RDATA_IM0(15) => RDATA_IM0(15), RDATA_IM0(14) => 
        RDATA_IM0(14), RDATA_IM0(13) => RDATA_IM0(13), 
        RDATA_IM0(12) => RDATA_IM0(12), RDATA_IM0(11) => 
        RDATA_IM0(11), RDATA_IM0(10) => RDATA_IM0(10), 
        RDATA_IM0(9) => RDATA_IM0(9), RDATA_IM0(8) => 
        RDATA_IM0(8), RDATA_IM0(7) => RDATA_IM0(7), RDATA_IM0(6)
         => RDATA_IM0(6), RDATA_IM0(5) => RDATA_IM0(5), 
        RDATA_IM0(4) => RDATA_IM0(4), RDATA_IM0(3) => 
        RDATA_IM0(3), RDATA_IM0(2) => RDATA_IM0(2), RDATA_IM0(1)
         => RDATA_IM0(1), RDATA_IM0(0) => RDATA_IM0(0), 
        axi_state_0 => axi_state_0, RDATA_reg_3 => RDATA_reg_3, 
        RDATA_reg_0 => RDATA_reg_0, COREAXI_0_AXImslave16_RDATA_3
         => COREAXI_0_AXImslave16_RDATA_3, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        COREAXI_0_AXImslave16_RDATA_0, 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        COREAXI_0_AXImslave16_RDATA_m_57, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        COREAXI_0_AXImslave16_RDATA_m_58, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        COREAXI_0_AXImslave16_RDATA_m_41, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        COREAXI_0_AXImslave16_RDATA_m_42, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        COREAXI_0_AXImslave16_RDATA_m_47, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        COREAXI_0_AXImslave16_RDATA_m_49, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        COREAXI_0_AXImslave16_RDATA_m_50, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        COREAXI_0_AXImslave16_RDATA_m_33, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        COREAXI_0_AXImslave16_RDATA_m_34, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        COREAXI_0_AXImslave16_RDATA_m_11, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        COREAXI_0_AXImslave16_RDATA_m_12, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        COREAXI_0_AXImslave16_RDATA_m_13, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        COREAXI_0_AXImslave16_RDATA_m_14, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        COREAXI_0_AXImslave16_RDATA_m_15, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        COREAXI_0_AXImslave16_RDATA_m_19, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        COREAXI_0_AXImslave16_RDATA_m_20, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        COREAXI_0_AXImslave16_RDATA_m_21, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        COREAXI_0_AXImslave16_RDATA_m_23, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        COREAXI_0_AXImslave16_RDATA_m_0, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        COREAXI_0_AXImslave16_RDATA_m_1, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        COREAXI_0_AXImslave16_RDATA_m_4, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        COREAXI_0_AXImslave16_RDATA_m_5, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        COREAXI_0_AXImslave16_RDATA_m_6, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        COREAXI_0_AXImslave16_RDATA_m_7, 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        COREAXI_0_AXImslave16_RDATA_m_8, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        COREAXI_0_AXImslave16_RDATA_m_9, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        COREAXI_0_AXImslave16_RDATA_m_10, BVALID_IM0 => 
        BVALID_IM0, COREAXI_0_AXImslave16_BVALID => 
        COREAXI_0_AXImslave16_BVALID, N_3297 => N_3297, 
        RREADY_MI0 => RREADY_MI0, N_389 => N_389, N_74 => N_74, 
        N_3167_i => N_3167_i, N_23 => N_23, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, RVALID_IM0 => 
        RVALID_IM0, RLAST_IM0 => RLAST_IM0, N_3170_i => N_3170_i, 
        N_39 => N_39, N_78_mux_i => N_78_mux_i, N_79_mux_i => 
        N_79_mux_i, N_80_mux_i => N_80_mux_i, N_70_mux_i => 
        N_70_mux_i, N_71_mux_i => N_71_mux_i, N_72_mux_i => 
        N_72_mux_i, N_3094_i => N_3094_i, N_3096_i => N_3096_i, 
        N_3098_i => N_3098_i, N_3100_i => N_3100_i, N_3102_i => 
        N_3102_i, N_3169_i => N_3169_i, N_3066_i => N_3066_i, 
        N_67_mux_i => N_67_mux_i, N_68_mux_i => N_68_mux_i, 
        N_69_mux_i => N_69_mux_i, N_75_mux_i => N_75_mux_i, 
        N_76_mux_i => N_76_mux_i, N_77_mux_i => N_77_mux_i, 
        i22_mux_2_i => i22_mux_2_i, i22_mux_3_i => i22_mux_3_i, 
        i22_mux_4_i => i22_mux_4_i, i22_mux_5_i => i22_mux_5_i, 
        N_8_i => N_8_i, i17_mux_2_i => i17_mux_2_i, N_3064_i => 
        N_3064_i, N_3092_i => N_3092_i, i17_mux_i => i17_mux_i, 
        i17_mux_0_i => i17_mux_0_i, i17_mux_1_i => i17_mux_1_i, 
        i22_mux_i => i22_mux_i, i22_mux_0_i => i22_mux_0_i, 
        i22_mux_1_i => i22_mux_1_i, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    WVALID_IS16_gated_r : SLE
      port map(D => WVALID_IS16_gated, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \WVALID_IS16_gated_r\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \AWVALID_IS16\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => \AWADDR_IS16_gated_r[27]_net_1\, B => 
        \AWVALID_IS16_gated_r\, C => AWVALID_IS16_gated, D => 
        \AWADDR_IS16_gated_r[26]_net_1\, Y => AWVALID_IS16);
    
    \ARVALID_IS16\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => \ARADDR_IS16_gated_r[27]_net_1\, B => 
        \ARVALID_IS16_gated_r\, C => ARVALID_IS16_gated, D => 
        \ARADDR_IS16_gated_r[26]_net_1\, Y => ARVALID_IS16);
    
    \ARADDR_IS16_gated_r[27]\ : SLE
      port map(D => \ARADDR_IS16_gated[27]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ARADDR_IS16_gated_r[27]_net_1\);
    
    \WVALID_IS16\ : CFG4
      generic map(INIT => x"40C0")

      port map(A => \AWADDR_IS16_gated_r[27]_net_1\, B => 
        \WVALID_IS16_gated_r\, C => WVALID_IS16_gated, D => 
        \AWADDR_IS16_gated_r[26]_net_1\, Y => WVALID_IS16);
    
    AWVALID_IS16_gated_r : SLE
      port map(D => AWVALID_IS16_gated, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWVALID_IS16_gated_r\);
    
    \AWADDR_IS16_gated_r[27]\ : SLE
      port map(D => \AWADDR_IS16_gated[27]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AWADDR_IS16_gated_r[27]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top_sb_COREAXI_0_COREAXI is

    port( COREAXI_0_AXImslave16_AWSIZE         : out   std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_ARADDR         : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_AWADDR         : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_WSTRB          : out   std_logic_vector(7 downto 0);
          COREAXI_0_AXImslave16_WDATA          : out   std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_ARSIZE         : out   std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : out   std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : in    std_logic_vector(63 downto 16);
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : in    std_logic_vector(27 downto 1);
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : in    std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_ARBURST_0      : out   std_logic;
          axi_current_state_0                  : in    std_logic;
          axi_current_state_3                  : in    std_logic;
          axi_state_0                          : in    std_logic;
          RDATA_reg_3                          : in    std_logic;
          RDATA_reg_0                          : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_3        : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_0        : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23     : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_8      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9      : in    std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10     : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic;
          COREAXI_0_AXImslave16_WVALID         : out   std_logic;
          WREADY_SI16_i                        : in    std_logic;
          COREAXI_0_AXImslave16_AWVALID        : out   std_logic;
          COREAXI_0_AXImslave16_AWREADY        : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : out   std_logic;
          wready_m_xhdl2                       : out   std_logic;
          N_1445_i                             : in    std_logic;
          N_1446_i                             : in    std_logic;
          N_1447_i                             : in    std_logic;
          N_1448_i                             : in    std_logic;
          N_1449_i                             : in    std_logic;
          N_1450_i                             : in    std_logic;
          N_1451_i                             : in    std_logic;
          N_1452_i                             : in    std_logic;
          N_202_i                              : in    std_logic;
          N_201_i                              : in    std_logic;
          N_200_i                              : in    std_logic;
          N_197_i                              : in    std_logic;
          N_195_i                              : in    std_logic;
          N_134_i                              : in    std_logic;
          N_133_i                              : in    std_logic;
          N_380_i                              : in    std_logic;
          N_278_i                              : in    std_logic;
          N_381_i                              : in    std_logic;
          N_382_i                              : in    std_logic;
          N_277_i                              : in    std_logic;
          N_276_i                              : in    std_logic;
          N_275_i                              : in    std_logic;
          N_274_i                              : in    std_logic;
          N_273_i                              : in    std_logic;
          N_272_i                              : in    std_logic;
          N_203_i                              : in    std_logic;
          N_137_i                              : in    std_logic;
          N_136_i                              : in    std_logic;
          N_135_i                              : in    std_logic;
          N_48                                 : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : out   std_logic;
          araddr_arvalid_clr_d                 : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : in    std_logic;
          awaddr_awvalid_clr_d                 : in    std_logic;
          MSS_READY                            : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          COREAXI_0_AXImslave16_BVALID         : in    std_logic;
          N_3297                               : in    std_logic;
          N_389                                : in    std_logic;
          N_74                                 : in    std_logic;
          N_3167_i                             : out   std_logic;
          N_23                                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic;
          N_3170_i                             : in    std_logic;
          N_39                                 : in    std_logic;
          N_78_mux_i                           : in    std_logic;
          N_79_mux_i                           : in    std_logic;
          N_80_mux_i                           : in    std_logic;
          N_70_mux_i                           : in    std_logic;
          N_71_mux_i                           : in    std_logic;
          N_72_mux_i                           : in    std_logic;
          N_3094_i                             : in    std_logic;
          N_3096_i                             : in    std_logic;
          N_3098_i                             : in    std_logic;
          N_3100_i                             : in    std_logic;
          N_3102_i                             : in    std_logic;
          N_3169_i                             : in    std_logic;
          N_3066_i                             : in    std_logic;
          N_67_mux_i                           : in    std_logic;
          N_68_mux_i                           : in    std_logic;
          N_69_mux_i                           : in    std_logic;
          N_75_mux_i                           : in    std_logic;
          N_76_mux_i                           : in    std_logic;
          N_77_mux_i                           : in    std_logic;
          i22_mux_2_i                          : in    std_logic;
          i22_mux_3_i                          : in    std_logic;
          i22_mux_4_i                          : in    std_logic;
          i22_mux_5_i                          : in    std_logic;
          N_8_i                                : in    std_logic;
          i17_mux_2_i                          : in    std_logic;
          N_3064_i                             : in    std_logic;
          N_3092_i                             : in    std_logic;
          i17_mux_i                            : in    std_logic;
          i17_mux_0_i                          : in    std_logic;
          i17_mux_1_i                          : in    std_logic;
          i22_mux_i                            : in    std_logic;
          i22_mux_0_i                          : in    std_logic;
          i22_mux_1_i                          : in    std_logic;
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic;
          COREAXI_0_AXImslave16_ARVALID        : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic;
          WREADY_SI16                          : in    std_logic;
          N_75_i                               : in    std_logic
        );

end top_sb_COREAXI_0_COREAXI;

architecture DEF_ARCH of top_sb_COREAXI_0_COREAXI is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component axi_slave_stage
    port( AWSIZE_IS16_gated               : in    std_logic_vector(1 downto 0) := (others => 'U');
          ARADDR_IS16_gated               : in    std_logic_vector(23 downto 1) := (others => 'U');
          AWADDR_IS16_gated               : in    std_logic_vector(23 downto 1) := (others => 'U');
          ARSIZE_IS16_gated               : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_ARSIZE    : out   std_logic_vector(1 downto 0);
          WDATA_IS16_gated                : in    std_logic_vector(63 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_WDATA     : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated                : in    std_logic_vector(7 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_WSTRB     : out   std_logic_vector(7 downto 0);
          COREAXI_0_AXImslave16_AWADDR    : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_ARADDR    : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_AWSIZE    : out   std_logic_vector(1 downto 0);
          ARBURST_IS16_gated_0            : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARBURST_0 : out   std_logic;
          WREADY_SI16                     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_AWREADY   : in    std_logic := 'U';
          WVALID_IS16                     : in    std_logic := 'U';
          AWVALID_IS16                    : in    std_logic := 'U';
          ARVALID_IS16                    : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID   : out   std_logic;
          AWREADY_SI16                    : out   std_logic;
          COREAXI_0_AXImslave16_AWVALID   : out   std_logic;
          WREADY_SI16_i                   : in    std_logic := 'U';
          COREAXI_0_AXImslave16_WVALID    : out   std_logic;
          SDRCLK_c                        : in    std_logic := 'U';
          MSS_READY                       : in    std_logic := 'U'
        );
  end component;

  component axi_master_stage
    port( RDATA_IM0                            : in    std_logic_vector(63 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : in    std_logic_vector(27 downto 1) := (others => 'U');
          AWADDR_MI0                           : out   std_logic_vector(27 downto 1);
          ARADDR_MI0                           : out   std_logic_vector(27 downto 1);
          ARSIZE_MI0                           : out   std_logic_vector(1 downto 0);
          AWSIZE_MI0                           : out   std_logic_vector(1 downto 0);
          WDATA_MI0                            : out   std_logic_vector(63 downto 0);
          WSTRB_MI0                            : out   std_logic_vector(7 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : in    std_logic_vector(63 downto 16) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : out   std_logic_vector(63 downto 0);
          axi_current_state_0                  : in    std_logic := 'U';
          axi_current_state_3                  : in    std_logic := 'U';
          ARBURST_MI0_0                        : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          AWLOCK_MI0_i_0                       : out   std_logic;
          ARLOCK_MI0_i_0                       : out   std_logic;
          ARREADY_IM0                          : in    std_logic := 'U';
          awaddr_awvalid_clr_d                 : in    std_logic := 'U';
          RVALID_IM0                           : in    std_logic := 'U';
          RLAST_IM0                            : in    std_logic := 'U';
          AWREADY_IM0                          : in    std_logic := 'U';
          WREADY_IM0                           : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : in    std_logic := 'U';
          RREADY_MI0                           : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic := 'U';
          araddr_arvalid_clr_d                 : in    std_logic := 'U';
          BVALID_IM0                           : in    std_logic := 'U';
          m0_rd_end                            : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : out   std_logic;
          m0_wr_end                            : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : out   std_logic;
          WVALID_MI0                           : out   std_logic;
          N_48                                 : in    std_logic := 'U';
          AWVALID_MI0                          : out   std_logic;
          ARVALID_MI0                          : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          N_75_i                               : in    std_logic := 'U';
          N_135_i                              : in    std_logic := 'U';
          N_136_i                              : in    std_logic := 'U';
          N_137_i                              : in    std_logic := 'U';
          N_203_i                              : in    std_logic := 'U';
          N_272_i                              : in    std_logic := 'U';
          N_273_i                              : in    std_logic := 'U';
          N_274_i                              : in    std_logic := 'U';
          N_275_i                              : in    std_logic := 'U';
          N_276_i                              : in    std_logic := 'U';
          N_277_i                              : in    std_logic := 'U';
          N_382_i                              : in    std_logic := 'U';
          N_381_i                              : in    std_logic := 'U';
          N_278_i                              : in    std_logic := 'U';
          N_380_i                              : in    std_logic := 'U';
          N_133_i                              : in    std_logic := 'U';
          N_134_i                              : in    std_logic := 'U';
          N_195_i                              : in    std_logic := 'U';
          N_197_i                              : in    std_logic := 'U';
          N_200_i                              : in    std_logic := 'U';
          N_201_i                              : in    std_logic := 'U';
          N_202_i                              : in    std_logic := 'U';
          N_1452_i                             : in    std_logic := 'U';
          N_1451_i                             : in    std_logic := 'U';
          N_1450_i                             : in    std_logic := 'U';
          N_1449_i                             : in    std_logic := 'U';
          N_1448_i                             : in    std_logic := 'U';
          N_1447_i                             : in    std_logic := 'U';
          N_1446_i                             : in    std_logic := 'U';
          N_1445_i                             : in    std_logic := 'U';
          wready_m_xhdl2                       : out   std_logic;
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : out   std_logic
        );
  end component;

  component axi_interconnect_ntom
    port( AWSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          AWADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          AWADDR_IS16_gated                    : out   std_logic_vector(23 downto 1);
          AWSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          WDATA_MI0                            : in    std_logic_vector(63 downto 0) := (others => 'U');
          WSTRB_MI0                            : in    std_logic_vector(7 downto 0) := (others => 'U');
          WDATA_IS16_gated                     : out   std_logic_vector(63 downto 0);
          WSTRB_IS16_gated                     : out   std_logic_vector(7 downto 0);
          ARSIZE_IS16_gated                    : out   std_logic_vector(1 downto 0);
          ARADDR_MI0                           : in    std_logic_vector(27 downto 1) := (others => 'U');
          ARADDR_IS16_gated                    : out   std_logic_vector(23 downto 1);
          ARSIZE_MI0                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          RDATA_IM0                            : out   std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          AWLOCK_MI0_i_0                       : in    std_logic := 'U';
          ARBURST_IS16_gated_0                 : out   std_logic;
          ARBURST_MI0_0                        : in    std_logic := 'U';
          ARLOCK_MI0_i_0                       : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_57     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_58     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_41     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_42     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_47     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_49     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_50     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_33     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_34     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_11     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_12     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_13     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_14     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_15     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_19     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_20     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_21     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_23     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_0      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_1      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_4      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_5      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_6      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_7      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_8      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_9      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_10     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_3        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_0        : in    std_logic := 'U';
          RDATA_reg_3                          : in    std_logic := 'U';
          RDATA_reg_0                          : in    std_logic := 'U';
          axi_state_0                          : in    std_logic := 'U';
          AWREADY_IM0                          : out   std_logic;
          N_75_i                               : in    std_logic := 'U';
          AWVALID_MI0                          : in    std_logic := 'U';
          AWREADY_SI16                         : in    std_logic := 'U';
          m0_wr_end                            : in    std_logic := 'U';
          WREADY_SI16                          : in    std_logic := 'U';
          WVALID_MI0                           : in    std_logic := 'U';
          WREADY_IM0                           : out   std_logic;
          ARREADY_IM0                          : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic := 'U';
          ARVALID_MI0                          : in    std_logic := 'U';
          m0_rd_end                            : in    std_logic := 'U';
          i22_mux_1_i                          : in    std_logic := 'U';
          i22_mux_0_i                          : in    std_logic := 'U';
          i22_mux_i                            : in    std_logic := 'U';
          i17_mux_1_i                          : in    std_logic := 'U';
          i17_mux_0_i                          : in    std_logic := 'U';
          i17_mux_i                            : in    std_logic := 'U';
          N_3092_i                             : in    std_logic := 'U';
          N_3064_i                             : in    std_logic := 'U';
          i17_mux_2_i                          : in    std_logic := 'U';
          N_8_i                                : in    std_logic := 'U';
          i22_mux_5_i                          : in    std_logic := 'U';
          i22_mux_4_i                          : in    std_logic := 'U';
          i22_mux_3_i                          : in    std_logic := 'U';
          i22_mux_2_i                          : in    std_logic := 'U';
          N_77_mux_i                           : in    std_logic := 'U';
          N_76_mux_i                           : in    std_logic := 'U';
          N_75_mux_i                           : in    std_logic := 'U';
          N_69_mux_i                           : in    std_logic := 'U';
          N_68_mux_i                           : in    std_logic := 'U';
          N_67_mux_i                           : in    std_logic := 'U';
          N_3066_i                             : in    std_logic := 'U';
          N_3169_i                             : in    std_logic := 'U';
          N_3102_i                             : in    std_logic := 'U';
          N_3100_i                             : in    std_logic := 'U';
          N_3098_i                             : in    std_logic := 'U';
          N_3096_i                             : in    std_logic := 'U';
          N_3094_i                             : in    std_logic := 'U';
          N_72_mux_i                           : in    std_logic := 'U';
          N_71_mux_i                           : in    std_logic := 'U';
          N_70_mux_i                           : in    std_logic := 'U';
          N_80_mux_i                           : in    std_logic := 'U';
          N_79_mux_i                           : in    std_logic := 'U';
          N_78_mux_i                           : in    std_logic := 'U';
          N_39                                 : in    std_logic := 'U';
          N_3170_i                             : in    std_logic := 'U';
          RLAST_IM0                            : out   std_logic;
          RVALID_IM0                           : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic := 'U';
          N_23                                 : out   std_logic;
          N_3167_i                             : out   std_logic;
          N_74                                 : in    std_logic := 'U';
          N_389                                : in    std_logic := 'U';
          RREADY_MI0                           : in    std_logic := 'U';
          N_3297                               : in    std_logic := 'U';
          COREAXI_0_AXImslave16_BVALID         : in    std_logic := 'U';
          BVALID_IM0                           : out   std_logic;
          ARVALID_IS16                         : out   std_logic;
          AWVALID_IS16                         : out   std_logic;
          WVALID_IS16                          : out   std_logic;
          SDRCLK_c                             : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \AWSIZE_IS16_gated[0]\, \AWSIZE_IS16_gated[1]\, 
        \AWADDR_MI0[1]\, \AWADDR_MI0[2]\, \AWADDR_MI0[3]\, 
        \AWADDR_MI0[4]\, \AWADDR_MI0[5]\, \AWADDR_MI0[6]\, 
        \AWADDR_MI0[7]\, \AWADDR_MI0[8]\, \AWADDR_MI0[9]\, 
        \AWADDR_MI0[10]\, \AWADDR_MI0[11]\, \AWADDR_MI0[12]\, 
        \AWADDR_MI0[13]\, \AWADDR_MI0[14]\, \AWADDR_MI0[15]\, 
        \AWADDR_MI0[16]\, \AWADDR_MI0[17]\, \AWADDR_MI0[18]\, 
        \AWADDR_MI0[19]\, \AWADDR_MI0[20]\, \AWADDR_MI0[21]\, 
        \AWADDR_MI0[22]\, \AWADDR_MI0[23]\, \AWADDR_MI0[26]\, 
        \AWADDR_MI0[27]\, \AWADDR_IS16_gated[1]\, 
        \AWADDR_IS16_gated[2]\, \AWADDR_IS16_gated[3]\, 
        \AWADDR_IS16_gated[4]\, \AWADDR_IS16_gated[5]\, 
        \AWADDR_IS16_gated[6]\, \AWADDR_IS16_gated[7]\, 
        \AWADDR_IS16_gated[8]\, \AWADDR_IS16_gated[9]\, 
        \AWADDR_IS16_gated[10]\, \AWADDR_IS16_gated[11]\, 
        \AWADDR_IS16_gated[12]\, \AWADDR_IS16_gated[13]\, 
        \AWADDR_IS16_gated[14]\, \AWADDR_IS16_gated[15]\, 
        \AWADDR_IS16_gated[16]\, \AWADDR_IS16_gated[17]\, 
        \AWADDR_IS16_gated[18]\, \AWADDR_IS16_gated[19]\, 
        \AWADDR_IS16_gated[20]\, \AWADDR_IS16_gated[21]\, 
        \AWADDR_IS16_gated[22]\, \AWADDR_IS16_gated[23]\, 
        \AWSIZE_MI0[0]\, \AWSIZE_MI0[1]\, \AWLOCK_MI0_i[1]\, 
        \WDATA_MI0[0]\, \WDATA_MI0[1]\, \WDATA_MI0[2]\, 
        \WDATA_MI0[3]\, \WDATA_MI0[4]\, \WDATA_MI0[5]\, 
        \WDATA_MI0[6]\, \WDATA_MI0[7]\, \WDATA_MI0[8]\, 
        \WDATA_MI0[9]\, \WDATA_MI0[10]\, \WDATA_MI0[11]\, 
        \WDATA_MI0[12]\, \WDATA_MI0[13]\, \WDATA_MI0[14]\, 
        \WDATA_MI0[15]\, \WDATA_MI0[16]\, \WDATA_MI0[17]\, 
        \WDATA_MI0[18]\, \WDATA_MI0[19]\, \WDATA_MI0[20]\, 
        \WDATA_MI0[21]\, \WDATA_MI0[22]\, \WDATA_MI0[23]\, 
        \WDATA_MI0[24]\, \WDATA_MI0[25]\, \WDATA_MI0[26]\, 
        \WDATA_MI0[27]\, \WDATA_MI0[28]\, \WDATA_MI0[29]\, 
        \WDATA_MI0[30]\, \WDATA_MI0[31]\, \WDATA_MI0[32]\, 
        \WDATA_MI0[33]\, \WDATA_MI0[34]\, \WDATA_MI0[35]\, 
        \WDATA_MI0[36]\, \WDATA_MI0[37]\, \WDATA_MI0[38]\, 
        \WDATA_MI0[39]\, \WDATA_MI0[40]\, \WDATA_MI0[41]\, 
        \WDATA_MI0[42]\, \WDATA_MI0[43]\, \WDATA_MI0[44]\, 
        \WDATA_MI0[45]\, \WDATA_MI0[46]\, \WDATA_MI0[47]\, 
        \WDATA_MI0[48]\, \WDATA_MI0[49]\, \WDATA_MI0[50]\, 
        \WDATA_MI0[51]\, \WDATA_MI0[52]\, \WDATA_MI0[53]\, 
        \WDATA_MI0[54]\, \WDATA_MI0[55]\, \WDATA_MI0[56]\, 
        \WDATA_MI0[57]\, \WDATA_MI0[58]\, \WDATA_MI0[59]\, 
        \WDATA_MI0[60]\, \WDATA_MI0[61]\, \WDATA_MI0[62]\, 
        \WDATA_MI0[63]\, \WSTRB_MI0[0]\, \WSTRB_MI0[1]\, 
        \WSTRB_MI0[2]\, \WSTRB_MI0[3]\, \WSTRB_MI0[4]\, 
        \WSTRB_MI0[5]\, \WSTRB_MI0[6]\, \WSTRB_MI0[7]\, 
        \WDATA_IS16_gated[0]\, \WDATA_IS16_gated[1]\, 
        \WDATA_IS16_gated[2]\, \WDATA_IS16_gated[3]\, 
        \WDATA_IS16_gated[4]\, \WDATA_IS16_gated[5]\, 
        \WDATA_IS16_gated[6]\, \WDATA_IS16_gated[7]\, 
        \WDATA_IS16_gated[8]\, \WDATA_IS16_gated[9]\, 
        \WDATA_IS16_gated[10]\, \WDATA_IS16_gated[11]\, 
        \WDATA_IS16_gated[12]\, \WDATA_IS16_gated[13]\, 
        \WDATA_IS16_gated[14]\, \WDATA_IS16_gated[15]\, 
        \WDATA_IS16_gated[16]\, \WDATA_IS16_gated[17]\, 
        \WDATA_IS16_gated[18]\, \WDATA_IS16_gated[19]\, 
        \WDATA_IS16_gated[20]\, \WDATA_IS16_gated[21]\, 
        \WDATA_IS16_gated[22]\, \WDATA_IS16_gated[23]\, 
        \WDATA_IS16_gated[24]\, \WDATA_IS16_gated[25]\, 
        \WDATA_IS16_gated[26]\, \WDATA_IS16_gated[27]\, 
        \WDATA_IS16_gated[28]\, \WDATA_IS16_gated[29]\, 
        \WDATA_IS16_gated[30]\, \WDATA_IS16_gated[31]\, 
        \WDATA_IS16_gated[32]\, \WDATA_IS16_gated[33]\, 
        \WDATA_IS16_gated[34]\, \WDATA_IS16_gated[35]\, 
        \WDATA_IS16_gated[36]\, \WDATA_IS16_gated[37]\, 
        \WDATA_IS16_gated[38]\, \WDATA_IS16_gated[39]\, 
        \WDATA_IS16_gated[40]\, \WDATA_IS16_gated[41]\, 
        \WDATA_IS16_gated[42]\, \WDATA_IS16_gated[43]\, 
        \WDATA_IS16_gated[44]\, \WDATA_IS16_gated[45]\, 
        \WDATA_IS16_gated[46]\, \WDATA_IS16_gated[47]\, 
        \WDATA_IS16_gated[48]\, \WDATA_IS16_gated[49]\, 
        \WDATA_IS16_gated[50]\, \WDATA_IS16_gated[51]\, 
        \WDATA_IS16_gated[52]\, \WDATA_IS16_gated[53]\, 
        \WDATA_IS16_gated[54]\, \WDATA_IS16_gated[55]\, 
        \WDATA_IS16_gated[56]\, \WDATA_IS16_gated[57]\, 
        \WDATA_IS16_gated[58]\, \WDATA_IS16_gated[59]\, 
        \WDATA_IS16_gated[60]\, \WDATA_IS16_gated[61]\, 
        \WDATA_IS16_gated[62]\, \WDATA_IS16_gated[63]\, 
        \WSTRB_IS16_gated[0]\, \WSTRB_IS16_gated[1]\, 
        \WSTRB_IS16_gated[2]\, \WSTRB_IS16_gated[3]\, 
        \WSTRB_IS16_gated[4]\, \WSTRB_IS16_gated[5]\, 
        \WSTRB_IS16_gated[6]\, \WSTRB_IS16_gated[7]\, 
        \ARBURST_IS16_gated[0]\, \ARSIZE_IS16_gated[0]\, 
        \ARSIZE_IS16_gated[1]\, \ARADDR_MI0[1]\, \ARADDR_MI0[2]\, 
        \ARADDR_MI0[3]\, \ARADDR_MI0[4]\, \ARADDR_MI0[5]\, 
        \ARADDR_MI0[6]\, \ARADDR_MI0[7]\, \ARADDR_MI0[8]\, 
        \ARADDR_MI0[9]\, \ARADDR_MI0[10]\, \ARADDR_MI0[11]\, 
        \ARADDR_MI0[12]\, \ARADDR_MI0[13]\, \ARADDR_MI0[14]\, 
        \ARADDR_MI0[15]\, \ARADDR_MI0[16]\, \ARADDR_MI0[17]\, 
        \ARADDR_MI0[18]\, \ARADDR_MI0[19]\, \ARADDR_MI0[20]\, 
        \ARADDR_MI0[21]\, \ARADDR_MI0[22]\, \ARADDR_MI0[23]\, 
        \ARADDR_MI0[26]\, \ARADDR_MI0[27]\, 
        \ARADDR_IS16_gated[1]\, \ARADDR_IS16_gated[2]\, 
        \ARADDR_IS16_gated[3]\, \ARADDR_IS16_gated[4]\, 
        \ARADDR_IS16_gated[5]\, \ARADDR_IS16_gated[6]\, 
        \ARADDR_IS16_gated[7]\, \ARADDR_IS16_gated[8]\, 
        \ARADDR_IS16_gated[9]\, \ARADDR_IS16_gated[10]\, 
        \ARADDR_IS16_gated[11]\, \ARADDR_IS16_gated[12]\, 
        \ARADDR_IS16_gated[13]\, \ARADDR_IS16_gated[14]\, 
        \ARADDR_IS16_gated[15]\, \ARADDR_IS16_gated[16]\, 
        \ARADDR_IS16_gated[17]\, \ARADDR_IS16_gated[18]\, 
        \ARADDR_IS16_gated[19]\, \ARADDR_IS16_gated[20]\, 
        \ARADDR_IS16_gated[21]\, \ARADDR_IS16_gated[22]\, 
        \ARADDR_IS16_gated[23]\, \ARBURST_MI0[0]\, 
        \ARSIZE_MI0[0]\, \ARSIZE_MI0[1]\, \ARLOCK_MI0_i[1]\, 
        \RDATA_IM0[0]\, \RDATA_IM0[1]\, \RDATA_IM0[2]\, 
        \RDATA_IM0[3]\, \RDATA_IM0[4]\, \RDATA_IM0[5]\, 
        \RDATA_IM0[6]\, \RDATA_IM0[7]\, \RDATA_IM0[8]\, 
        \RDATA_IM0[9]\, \RDATA_IM0[10]\, \RDATA_IM0[11]\, 
        \RDATA_IM0[12]\, \RDATA_IM0[13]\, \RDATA_IM0[14]\, 
        \RDATA_IM0[15]\, \RDATA_IM0[16]\, \RDATA_IM0[17]\, 
        \RDATA_IM0[18]\, \RDATA_IM0[19]\, \RDATA_IM0[20]\, 
        \RDATA_IM0[21]\, \RDATA_IM0[22]\, \RDATA_IM0[23]\, 
        \RDATA_IM0[24]\, \RDATA_IM0[25]\, \RDATA_IM0[26]\, 
        \RDATA_IM0[27]\, \RDATA_IM0[28]\, \RDATA_IM0[29]\, 
        \RDATA_IM0[30]\, \RDATA_IM0[31]\, \RDATA_IM0[32]\, 
        \RDATA_IM0[33]\, \RDATA_IM0[34]\, \RDATA_IM0[35]\, 
        \RDATA_IM0[36]\, \RDATA_IM0[37]\, \RDATA_IM0[38]\, 
        \RDATA_IM0[39]\, \RDATA_IM0[40]\, \RDATA_IM0[41]\, 
        \RDATA_IM0[42]\, \RDATA_IM0[43]\, \RDATA_IM0[44]\, 
        \RDATA_IM0[45]\, \RDATA_IM0[46]\, \RDATA_IM0[47]\, 
        \RDATA_IM0[48]\, \RDATA_IM0[49]\, \RDATA_IM0[50]\, 
        \RDATA_IM0[51]\, \RDATA_IM0[52]\, \RDATA_IM0[53]\, 
        \RDATA_IM0[54]\, \RDATA_IM0[55]\, \RDATA_IM0[56]\, 
        \RDATA_IM0[57]\, \RDATA_IM0[58]\, \RDATA_IM0[59]\, 
        \RDATA_IM0[60]\, \RDATA_IM0[61]\, \RDATA_IM0[62]\, 
        \RDATA_IM0[63]\, AWREADY_IM0, AWVALID_MI0, AWREADY_SI16, 
        m0_wr_end, WVALID_MI0, WREADY_IM0, ARREADY_IM0, 
        \COREAXI_0_AXImslave16_ARVALID\, ARVALID_MI0, m0_rd_end, 
        RLAST_IM0, RVALID_IM0, 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\, RREADY_MI0, 
        BVALID_IM0, ARVALID_IS16, AWVALID_IS16, WVALID_IS16, 
        GND_net_1, VCC_net_1 : std_logic;
    signal nc7, nc6, nc12, nc5, nc1, nc9, nc13, nc8, nc4, nc11, 
        nc3, nc10, nc2 : std_logic;

    for all : axi_slave_stage
	Use entity work.axi_slave_stage(DEF_ARCH);
    for all : axi_master_stage
	Use entity work.axi_master_stage(DEF_ARCH);
    for all : axi_interconnect_ntom
	Use entity work.axi_interconnect_ntom(DEF_ARCH);
begin 

    COREAHBLTOAXI_0_AXIMasterIF_RVALID <= 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\;
    COREAXI_0_AXImslave16_ARVALID <= 
        \COREAXI_0_AXImslave16_ARVALID\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \L23.slave_stage16\ : axi_slave_stage
      port map(AWSIZE_IS16_gated(1) => \AWSIZE_IS16_gated[1]\, 
        AWSIZE_IS16_gated(0) => \AWSIZE_IS16_gated[0]\, 
        ARADDR_IS16_gated(23) => \ARADDR_IS16_gated[23]\, 
        ARADDR_IS16_gated(22) => \ARADDR_IS16_gated[22]\, 
        ARADDR_IS16_gated(21) => \ARADDR_IS16_gated[21]\, 
        ARADDR_IS16_gated(20) => \ARADDR_IS16_gated[20]\, 
        ARADDR_IS16_gated(19) => \ARADDR_IS16_gated[19]\, 
        ARADDR_IS16_gated(18) => \ARADDR_IS16_gated[18]\, 
        ARADDR_IS16_gated(17) => \ARADDR_IS16_gated[17]\, 
        ARADDR_IS16_gated(16) => \ARADDR_IS16_gated[16]\, 
        ARADDR_IS16_gated(15) => \ARADDR_IS16_gated[15]\, 
        ARADDR_IS16_gated(14) => \ARADDR_IS16_gated[14]\, 
        ARADDR_IS16_gated(13) => \ARADDR_IS16_gated[13]\, 
        ARADDR_IS16_gated(12) => \ARADDR_IS16_gated[12]\, 
        ARADDR_IS16_gated(11) => \ARADDR_IS16_gated[11]\, 
        ARADDR_IS16_gated(10) => \ARADDR_IS16_gated[10]\, 
        ARADDR_IS16_gated(9) => \ARADDR_IS16_gated[9]\, 
        ARADDR_IS16_gated(8) => \ARADDR_IS16_gated[8]\, 
        ARADDR_IS16_gated(7) => \ARADDR_IS16_gated[7]\, 
        ARADDR_IS16_gated(6) => \ARADDR_IS16_gated[6]\, 
        ARADDR_IS16_gated(5) => \ARADDR_IS16_gated[5]\, 
        ARADDR_IS16_gated(4) => \ARADDR_IS16_gated[4]\, 
        ARADDR_IS16_gated(3) => \ARADDR_IS16_gated[3]\, 
        ARADDR_IS16_gated(2) => \ARADDR_IS16_gated[2]\, 
        ARADDR_IS16_gated(1) => \ARADDR_IS16_gated[1]\, 
        AWADDR_IS16_gated(23) => \AWADDR_IS16_gated[23]\, 
        AWADDR_IS16_gated(22) => \AWADDR_IS16_gated[22]\, 
        AWADDR_IS16_gated(21) => \AWADDR_IS16_gated[21]\, 
        AWADDR_IS16_gated(20) => \AWADDR_IS16_gated[20]\, 
        AWADDR_IS16_gated(19) => \AWADDR_IS16_gated[19]\, 
        AWADDR_IS16_gated(18) => \AWADDR_IS16_gated[18]\, 
        AWADDR_IS16_gated(17) => \AWADDR_IS16_gated[17]\, 
        AWADDR_IS16_gated(16) => \AWADDR_IS16_gated[16]\, 
        AWADDR_IS16_gated(15) => \AWADDR_IS16_gated[15]\, 
        AWADDR_IS16_gated(14) => \AWADDR_IS16_gated[14]\, 
        AWADDR_IS16_gated(13) => \AWADDR_IS16_gated[13]\, 
        AWADDR_IS16_gated(12) => \AWADDR_IS16_gated[12]\, 
        AWADDR_IS16_gated(11) => \AWADDR_IS16_gated[11]\, 
        AWADDR_IS16_gated(10) => \AWADDR_IS16_gated[10]\, 
        AWADDR_IS16_gated(9) => \AWADDR_IS16_gated[9]\, 
        AWADDR_IS16_gated(8) => \AWADDR_IS16_gated[8]\, 
        AWADDR_IS16_gated(7) => \AWADDR_IS16_gated[7]\, 
        AWADDR_IS16_gated(6) => \AWADDR_IS16_gated[6]\, 
        AWADDR_IS16_gated(5) => \AWADDR_IS16_gated[5]\, 
        AWADDR_IS16_gated(4) => \AWADDR_IS16_gated[4]\, 
        AWADDR_IS16_gated(3) => \AWADDR_IS16_gated[3]\, 
        AWADDR_IS16_gated(2) => \AWADDR_IS16_gated[2]\, 
        AWADDR_IS16_gated(1) => \AWADDR_IS16_gated[1]\, 
        ARSIZE_IS16_gated(1) => \ARSIZE_IS16_gated[1]\, 
        ARSIZE_IS16_gated(0) => \ARSIZE_IS16_gated[0]\, 
        COREAXI_0_AXImslave16_ARSIZE(1) => 
        COREAXI_0_AXImslave16_ARSIZE(1), 
        COREAXI_0_AXImslave16_ARSIZE(0) => 
        COREAXI_0_AXImslave16_ARSIZE(0), WDATA_IS16_gated(63) => 
        \WDATA_IS16_gated[63]\, WDATA_IS16_gated(62) => 
        \WDATA_IS16_gated[62]\, WDATA_IS16_gated(61) => 
        \WDATA_IS16_gated[61]\, WDATA_IS16_gated(60) => 
        \WDATA_IS16_gated[60]\, WDATA_IS16_gated(59) => 
        \WDATA_IS16_gated[59]\, WDATA_IS16_gated(58) => 
        \WDATA_IS16_gated[58]\, WDATA_IS16_gated(57) => 
        \WDATA_IS16_gated[57]\, WDATA_IS16_gated(56) => 
        \WDATA_IS16_gated[56]\, WDATA_IS16_gated(55) => 
        \WDATA_IS16_gated[55]\, WDATA_IS16_gated(54) => 
        \WDATA_IS16_gated[54]\, WDATA_IS16_gated(53) => 
        \WDATA_IS16_gated[53]\, WDATA_IS16_gated(52) => 
        \WDATA_IS16_gated[52]\, WDATA_IS16_gated(51) => 
        \WDATA_IS16_gated[51]\, WDATA_IS16_gated(50) => 
        \WDATA_IS16_gated[50]\, WDATA_IS16_gated(49) => 
        \WDATA_IS16_gated[49]\, WDATA_IS16_gated(48) => 
        \WDATA_IS16_gated[48]\, WDATA_IS16_gated(47) => 
        \WDATA_IS16_gated[47]\, WDATA_IS16_gated(46) => 
        \WDATA_IS16_gated[46]\, WDATA_IS16_gated(45) => 
        \WDATA_IS16_gated[45]\, WDATA_IS16_gated(44) => 
        \WDATA_IS16_gated[44]\, WDATA_IS16_gated(43) => 
        \WDATA_IS16_gated[43]\, WDATA_IS16_gated(42) => 
        \WDATA_IS16_gated[42]\, WDATA_IS16_gated(41) => 
        \WDATA_IS16_gated[41]\, WDATA_IS16_gated(40) => 
        \WDATA_IS16_gated[40]\, WDATA_IS16_gated(39) => 
        \WDATA_IS16_gated[39]\, WDATA_IS16_gated(38) => 
        \WDATA_IS16_gated[38]\, WDATA_IS16_gated(37) => 
        \WDATA_IS16_gated[37]\, WDATA_IS16_gated(36) => 
        \WDATA_IS16_gated[36]\, WDATA_IS16_gated(35) => 
        \WDATA_IS16_gated[35]\, WDATA_IS16_gated(34) => 
        \WDATA_IS16_gated[34]\, WDATA_IS16_gated(33) => 
        \WDATA_IS16_gated[33]\, WDATA_IS16_gated(32) => 
        \WDATA_IS16_gated[32]\, WDATA_IS16_gated(31) => 
        \WDATA_IS16_gated[31]\, WDATA_IS16_gated(30) => 
        \WDATA_IS16_gated[30]\, WDATA_IS16_gated(29) => 
        \WDATA_IS16_gated[29]\, WDATA_IS16_gated(28) => 
        \WDATA_IS16_gated[28]\, WDATA_IS16_gated(27) => 
        \WDATA_IS16_gated[27]\, WDATA_IS16_gated(26) => 
        \WDATA_IS16_gated[26]\, WDATA_IS16_gated(25) => 
        \WDATA_IS16_gated[25]\, WDATA_IS16_gated(24) => 
        \WDATA_IS16_gated[24]\, WDATA_IS16_gated(23) => 
        \WDATA_IS16_gated[23]\, WDATA_IS16_gated(22) => 
        \WDATA_IS16_gated[22]\, WDATA_IS16_gated(21) => 
        \WDATA_IS16_gated[21]\, WDATA_IS16_gated(20) => 
        \WDATA_IS16_gated[20]\, WDATA_IS16_gated(19) => 
        \WDATA_IS16_gated[19]\, WDATA_IS16_gated(18) => 
        \WDATA_IS16_gated[18]\, WDATA_IS16_gated(17) => 
        \WDATA_IS16_gated[17]\, WDATA_IS16_gated(16) => 
        \WDATA_IS16_gated[16]\, WDATA_IS16_gated(15) => 
        \WDATA_IS16_gated[15]\, WDATA_IS16_gated(14) => 
        \WDATA_IS16_gated[14]\, WDATA_IS16_gated(13) => 
        \WDATA_IS16_gated[13]\, WDATA_IS16_gated(12) => 
        \WDATA_IS16_gated[12]\, WDATA_IS16_gated(11) => 
        \WDATA_IS16_gated[11]\, WDATA_IS16_gated(10) => 
        \WDATA_IS16_gated[10]\, WDATA_IS16_gated(9) => 
        \WDATA_IS16_gated[9]\, WDATA_IS16_gated(8) => 
        \WDATA_IS16_gated[8]\, WDATA_IS16_gated(7) => 
        \WDATA_IS16_gated[7]\, WDATA_IS16_gated(6) => 
        \WDATA_IS16_gated[6]\, WDATA_IS16_gated(5) => 
        \WDATA_IS16_gated[5]\, WDATA_IS16_gated(4) => 
        \WDATA_IS16_gated[4]\, WDATA_IS16_gated(3) => 
        \WDATA_IS16_gated[3]\, WDATA_IS16_gated(2) => 
        \WDATA_IS16_gated[2]\, WDATA_IS16_gated(1) => 
        \WDATA_IS16_gated[1]\, WDATA_IS16_gated(0) => 
        \WDATA_IS16_gated[0]\, COREAXI_0_AXImslave16_WDATA(63)
         => COREAXI_0_AXImslave16_WDATA(63), 
        COREAXI_0_AXImslave16_WDATA(62) => 
        COREAXI_0_AXImslave16_WDATA(62), 
        COREAXI_0_AXImslave16_WDATA(61) => 
        COREAXI_0_AXImslave16_WDATA(61), 
        COREAXI_0_AXImslave16_WDATA(60) => 
        COREAXI_0_AXImslave16_WDATA(60), 
        COREAXI_0_AXImslave16_WDATA(59) => 
        COREAXI_0_AXImslave16_WDATA(59), 
        COREAXI_0_AXImslave16_WDATA(58) => 
        COREAXI_0_AXImslave16_WDATA(58), 
        COREAXI_0_AXImslave16_WDATA(57) => 
        COREAXI_0_AXImslave16_WDATA(57), 
        COREAXI_0_AXImslave16_WDATA(56) => 
        COREAXI_0_AXImslave16_WDATA(56), 
        COREAXI_0_AXImslave16_WDATA(55) => 
        COREAXI_0_AXImslave16_WDATA(55), 
        COREAXI_0_AXImslave16_WDATA(54) => 
        COREAXI_0_AXImslave16_WDATA(54), 
        COREAXI_0_AXImslave16_WDATA(53) => 
        COREAXI_0_AXImslave16_WDATA(53), 
        COREAXI_0_AXImslave16_WDATA(52) => 
        COREAXI_0_AXImslave16_WDATA(52), 
        COREAXI_0_AXImslave16_WDATA(51) => 
        COREAXI_0_AXImslave16_WDATA(51), 
        COREAXI_0_AXImslave16_WDATA(50) => 
        COREAXI_0_AXImslave16_WDATA(50), 
        COREAXI_0_AXImslave16_WDATA(49) => 
        COREAXI_0_AXImslave16_WDATA(49), 
        COREAXI_0_AXImslave16_WDATA(48) => 
        COREAXI_0_AXImslave16_WDATA(48), 
        COREAXI_0_AXImslave16_WDATA(47) => 
        COREAXI_0_AXImslave16_WDATA(47), 
        COREAXI_0_AXImslave16_WDATA(46) => 
        COREAXI_0_AXImslave16_WDATA(46), 
        COREAXI_0_AXImslave16_WDATA(45) => 
        COREAXI_0_AXImslave16_WDATA(45), 
        COREAXI_0_AXImslave16_WDATA(44) => 
        COREAXI_0_AXImslave16_WDATA(44), 
        COREAXI_0_AXImslave16_WDATA(43) => 
        COREAXI_0_AXImslave16_WDATA(43), 
        COREAXI_0_AXImslave16_WDATA(42) => 
        COREAXI_0_AXImslave16_WDATA(42), 
        COREAXI_0_AXImslave16_WDATA(41) => 
        COREAXI_0_AXImslave16_WDATA(41), 
        COREAXI_0_AXImslave16_WDATA(40) => 
        COREAXI_0_AXImslave16_WDATA(40), 
        COREAXI_0_AXImslave16_WDATA(39) => 
        COREAXI_0_AXImslave16_WDATA(39), 
        COREAXI_0_AXImslave16_WDATA(38) => 
        COREAXI_0_AXImslave16_WDATA(38), 
        COREAXI_0_AXImslave16_WDATA(37) => 
        COREAXI_0_AXImslave16_WDATA(37), 
        COREAXI_0_AXImslave16_WDATA(36) => 
        COREAXI_0_AXImslave16_WDATA(36), 
        COREAXI_0_AXImslave16_WDATA(35) => 
        COREAXI_0_AXImslave16_WDATA(35), 
        COREAXI_0_AXImslave16_WDATA(34) => 
        COREAXI_0_AXImslave16_WDATA(34), 
        COREAXI_0_AXImslave16_WDATA(33) => 
        COREAXI_0_AXImslave16_WDATA(33), 
        COREAXI_0_AXImslave16_WDATA(32) => 
        COREAXI_0_AXImslave16_WDATA(32), 
        COREAXI_0_AXImslave16_WDATA(31) => 
        COREAXI_0_AXImslave16_WDATA(31), 
        COREAXI_0_AXImslave16_WDATA(30) => 
        COREAXI_0_AXImslave16_WDATA(30), 
        COREAXI_0_AXImslave16_WDATA(29) => 
        COREAXI_0_AXImslave16_WDATA(29), 
        COREAXI_0_AXImslave16_WDATA(28) => 
        COREAXI_0_AXImslave16_WDATA(28), 
        COREAXI_0_AXImslave16_WDATA(27) => 
        COREAXI_0_AXImslave16_WDATA(27), 
        COREAXI_0_AXImslave16_WDATA(26) => 
        COREAXI_0_AXImslave16_WDATA(26), 
        COREAXI_0_AXImslave16_WDATA(25) => 
        COREAXI_0_AXImslave16_WDATA(25), 
        COREAXI_0_AXImslave16_WDATA(24) => 
        COREAXI_0_AXImslave16_WDATA(24), 
        COREAXI_0_AXImslave16_WDATA(23) => 
        COREAXI_0_AXImslave16_WDATA(23), 
        COREAXI_0_AXImslave16_WDATA(22) => 
        COREAXI_0_AXImslave16_WDATA(22), 
        COREAXI_0_AXImslave16_WDATA(21) => 
        COREAXI_0_AXImslave16_WDATA(21), 
        COREAXI_0_AXImslave16_WDATA(20) => 
        COREAXI_0_AXImslave16_WDATA(20), 
        COREAXI_0_AXImslave16_WDATA(19) => 
        COREAXI_0_AXImslave16_WDATA(19), 
        COREAXI_0_AXImslave16_WDATA(18) => 
        COREAXI_0_AXImslave16_WDATA(18), 
        COREAXI_0_AXImslave16_WDATA(17) => 
        COREAXI_0_AXImslave16_WDATA(17), 
        COREAXI_0_AXImslave16_WDATA(16) => 
        COREAXI_0_AXImslave16_WDATA(16), 
        COREAXI_0_AXImslave16_WDATA(15) => 
        COREAXI_0_AXImslave16_WDATA(15), 
        COREAXI_0_AXImslave16_WDATA(14) => 
        COREAXI_0_AXImslave16_WDATA(14), 
        COREAXI_0_AXImslave16_WDATA(13) => 
        COREAXI_0_AXImslave16_WDATA(13), 
        COREAXI_0_AXImslave16_WDATA(12) => 
        COREAXI_0_AXImslave16_WDATA(12), 
        COREAXI_0_AXImslave16_WDATA(11) => 
        COREAXI_0_AXImslave16_WDATA(11), 
        COREAXI_0_AXImslave16_WDATA(10) => 
        COREAXI_0_AXImslave16_WDATA(10), 
        COREAXI_0_AXImslave16_WDATA(9) => 
        COREAXI_0_AXImslave16_WDATA(9), 
        COREAXI_0_AXImslave16_WDATA(8) => 
        COREAXI_0_AXImslave16_WDATA(8), 
        COREAXI_0_AXImslave16_WDATA(7) => 
        COREAXI_0_AXImslave16_WDATA(7), 
        COREAXI_0_AXImslave16_WDATA(6) => 
        COREAXI_0_AXImslave16_WDATA(6), 
        COREAXI_0_AXImslave16_WDATA(5) => 
        COREAXI_0_AXImslave16_WDATA(5), 
        COREAXI_0_AXImslave16_WDATA(4) => 
        COREAXI_0_AXImslave16_WDATA(4), 
        COREAXI_0_AXImslave16_WDATA(3) => 
        COREAXI_0_AXImslave16_WDATA(3), 
        COREAXI_0_AXImslave16_WDATA(2) => 
        COREAXI_0_AXImslave16_WDATA(2), 
        COREAXI_0_AXImslave16_WDATA(1) => 
        COREAXI_0_AXImslave16_WDATA(1), 
        COREAXI_0_AXImslave16_WDATA(0) => 
        COREAXI_0_AXImslave16_WDATA(0), WSTRB_IS16_gated(7) => 
        \WSTRB_IS16_gated[7]\, WSTRB_IS16_gated(6) => 
        \WSTRB_IS16_gated[6]\, WSTRB_IS16_gated(5) => 
        \WSTRB_IS16_gated[5]\, WSTRB_IS16_gated(4) => 
        \WSTRB_IS16_gated[4]\, WSTRB_IS16_gated(3) => 
        \WSTRB_IS16_gated[3]\, WSTRB_IS16_gated(2) => 
        \WSTRB_IS16_gated[2]\, WSTRB_IS16_gated(1) => 
        \WSTRB_IS16_gated[1]\, WSTRB_IS16_gated(0) => 
        \WSTRB_IS16_gated[0]\, COREAXI_0_AXImslave16_WSTRB(7) => 
        COREAXI_0_AXImslave16_WSTRB(7), 
        COREAXI_0_AXImslave16_WSTRB(6) => 
        COREAXI_0_AXImslave16_WSTRB(6), 
        COREAXI_0_AXImslave16_WSTRB(5) => 
        COREAXI_0_AXImslave16_WSTRB(5), 
        COREAXI_0_AXImslave16_WSTRB(4) => 
        COREAXI_0_AXImslave16_WSTRB(4), 
        COREAXI_0_AXImslave16_WSTRB(3) => 
        COREAXI_0_AXImslave16_WSTRB(3), 
        COREAXI_0_AXImslave16_WSTRB(2) => 
        COREAXI_0_AXImslave16_WSTRB(2), 
        COREAXI_0_AXImslave16_WSTRB(1) => 
        COREAXI_0_AXImslave16_WSTRB(1), 
        COREAXI_0_AXImslave16_WSTRB(0) => 
        COREAXI_0_AXImslave16_WSTRB(0), 
        COREAXI_0_AXImslave16_AWADDR(23) => 
        COREAXI_0_AXImslave16_AWADDR(23), 
        COREAXI_0_AXImslave16_AWADDR(22) => 
        COREAXI_0_AXImslave16_AWADDR(22), 
        COREAXI_0_AXImslave16_AWADDR(21) => 
        COREAXI_0_AXImslave16_AWADDR(21), 
        COREAXI_0_AXImslave16_AWADDR(20) => 
        COREAXI_0_AXImslave16_AWADDR(20), 
        COREAXI_0_AXImslave16_AWADDR(19) => 
        COREAXI_0_AXImslave16_AWADDR(19), 
        COREAXI_0_AXImslave16_AWADDR(18) => 
        COREAXI_0_AXImslave16_AWADDR(18), 
        COREAXI_0_AXImslave16_AWADDR(17) => 
        COREAXI_0_AXImslave16_AWADDR(17), 
        COREAXI_0_AXImslave16_AWADDR(16) => 
        COREAXI_0_AXImslave16_AWADDR(16), 
        COREAXI_0_AXImslave16_AWADDR(15) => 
        COREAXI_0_AXImslave16_AWADDR(15), 
        COREAXI_0_AXImslave16_AWADDR(14) => 
        COREAXI_0_AXImslave16_AWADDR(14), 
        COREAXI_0_AXImslave16_AWADDR(13) => 
        COREAXI_0_AXImslave16_AWADDR(13), 
        COREAXI_0_AXImslave16_AWADDR(12) => 
        COREAXI_0_AXImslave16_AWADDR(12), 
        COREAXI_0_AXImslave16_AWADDR(11) => 
        COREAXI_0_AXImslave16_AWADDR(11), 
        COREAXI_0_AXImslave16_AWADDR(10) => 
        COREAXI_0_AXImslave16_AWADDR(10), 
        COREAXI_0_AXImslave16_AWADDR(9) => 
        COREAXI_0_AXImslave16_AWADDR(9), 
        COREAXI_0_AXImslave16_AWADDR(8) => 
        COREAXI_0_AXImslave16_AWADDR(8), 
        COREAXI_0_AXImslave16_AWADDR(7) => 
        COREAXI_0_AXImslave16_AWADDR(7), 
        COREAXI_0_AXImslave16_AWADDR(6) => 
        COREAXI_0_AXImslave16_AWADDR(6), 
        COREAXI_0_AXImslave16_AWADDR(5) => 
        COREAXI_0_AXImslave16_AWADDR(5), 
        COREAXI_0_AXImslave16_AWADDR(4) => 
        COREAXI_0_AXImslave16_AWADDR(4), 
        COREAXI_0_AXImslave16_AWADDR(3) => 
        COREAXI_0_AXImslave16_AWADDR(3), 
        COREAXI_0_AXImslave16_AWADDR(2) => 
        COREAXI_0_AXImslave16_AWADDR(2), 
        COREAXI_0_AXImslave16_AWADDR(1) => 
        COREAXI_0_AXImslave16_AWADDR(1), 
        COREAXI_0_AXImslave16_ARADDR(23) => 
        COREAXI_0_AXImslave16_ARADDR(23), 
        COREAXI_0_AXImslave16_ARADDR(22) => 
        COREAXI_0_AXImslave16_ARADDR(22), 
        COREAXI_0_AXImslave16_ARADDR(21) => 
        COREAXI_0_AXImslave16_ARADDR(21), 
        COREAXI_0_AXImslave16_ARADDR(20) => 
        COREAXI_0_AXImslave16_ARADDR(20), 
        COREAXI_0_AXImslave16_ARADDR(19) => 
        COREAXI_0_AXImslave16_ARADDR(19), 
        COREAXI_0_AXImslave16_ARADDR(18) => 
        COREAXI_0_AXImslave16_ARADDR(18), 
        COREAXI_0_AXImslave16_ARADDR(17) => 
        COREAXI_0_AXImslave16_ARADDR(17), 
        COREAXI_0_AXImslave16_ARADDR(16) => 
        COREAXI_0_AXImslave16_ARADDR(16), 
        COREAXI_0_AXImslave16_ARADDR(15) => 
        COREAXI_0_AXImslave16_ARADDR(15), 
        COREAXI_0_AXImslave16_ARADDR(14) => 
        COREAXI_0_AXImslave16_ARADDR(14), 
        COREAXI_0_AXImslave16_ARADDR(13) => 
        COREAXI_0_AXImslave16_ARADDR(13), 
        COREAXI_0_AXImslave16_ARADDR(12) => 
        COREAXI_0_AXImslave16_ARADDR(12), 
        COREAXI_0_AXImslave16_ARADDR(11) => 
        COREAXI_0_AXImslave16_ARADDR(11), 
        COREAXI_0_AXImslave16_ARADDR(10) => 
        COREAXI_0_AXImslave16_ARADDR(10), 
        COREAXI_0_AXImslave16_ARADDR(9) => 
        COREAXI_0_AXImslave16_ARADDR(9), 
        COREAXI_0_AXImslave16_ARADDR(8) => 
        COREAXI_0_AXImslave16_ARADDR(8), 
        COREAXI_0_AXImslave16_ARADDR(7) => 
        COREAXI_0_AXImslave16_ARADDR(7), 
        COREAXI_0_AXImslave16_ARADDR(6) => 
        COREAXI_0_AXImslave16_ARADDR(6), 
        COREAXI_0_AXImslave16_ARADDR(5) => 
        COREAXI_0_AXImslave16_ARADDR(5), 
        COREAXI_0_AXImslave16_ARADDR(4) => 
        COREAXI_0_AXImslave16_ARADDR(4), 
        COREAXI_0_AXImslave16_ARADDR(3) => 
        COREAXI_0_AXImslave16_ARADDR(3), 
        COREAXI_0_AXImslave16_ARADDR(2) => 
        COREAXI_0_AXImslave16_ARADDR(2), 
        COREAXI_0_AXImslave16_ARADDR(1) => 
        COREAXI_0_AXImslave16_ARADDR(1), 
        COREAXI_0_AXImslave16_AWSIZE(1) => 
        COREAXI_0_AXImslave16_AWSIZE(1), 
        COREAXI_0_AXImslave16_AWSIZE(0) => 
        COREAXI_0_AXImslave16_AWSIZE(0), ARBURST_IS16_gated_0 => 
        \ARBURST_IS16_gated[0]\, COREAXI_0_AXImslave16_ARBURST_0
         => COREAXI_0_AXImslave16_ARBURST_0, WREADY_SI16 => 
        WREADY_SI16, COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, 
        COREAXI_0_AXImslave16_AWREADY => 
        COREAXI_0_AXImslave16_AWREADY, WVALID_IS16 => WVALID_IS16, 
        AWVALID_IS16 => AWVALID_IS16, ARVALID_IS16 => 
        ARVALID_IS16, COREAXI_0_AXImslave16_ARVALID => 
        \COREAXI_0_AXImslave16_ARVALID\, AWREADY_SI16 => 
        AWREADY_SI16, COREAXI_0_AXImslave16_AWVALID => 
        COREAXI_0_AXImslave16_AWVALID, WREADY_SI16_i => 
        WREADY_SI16_i, COREAXI_0_AXImslave16_WVALID => 
        COREAXI_0_AXImslave16_WVALID, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY);
    
    \L3.master_stage0\ : axi_master_stage
      port map(RDATA_IM0(63) => \RDATA_IM0[63]\, RDATA_IM0(62)
         => \RDATA_IM0[62]\, RDATA_IM0(61) => \RDATA_IM0[61]\, 
        RDATA_IM0(60) => \RDATA_IM0[60]\, RDATA_IM0(59) => 
        \RDATA_IM0[59]\, RDATA_IM0(58) => \RDATA_IM0[58]\, 
        RDATA_IM0(57) => \RDATA_IM0[57]\, RDATA_IM0(56) => 
        \RDATA_IM0[56]\, RDATA_IM0(55) => \RDATA_IM0[55]\, 
        RDATA_IM0(54) => \RDATA_IM0[54]\, RDATA_IM0(53) => 
        \RDATA_IM0[53]\, RDATA_IM0(52) => \RDATA_IM0[52]\, 
        RDATA_IM0(51) => \RDATA_IM0[51]\, RDATA_IM0(50) => 
        \RDATA_IM0[50]\, RDATA_IM0(49) => \RDATA_IM0[49]\, 
        RDATA_IM0(48) => \RDATA_IM0[48]\, RDATA_IM0(47) => 
        \RDATA_IM0[47]\, RDATA_IM0(46) => \RDATA_IM0[46]\, 
        RDATA_IM0(45) => \RDATA_IM0[45]\, RDATA_IM0(44) => 
        \RDATA_IM0[44]\, RDATA_IM0(43) => \RDATA_IM0[43]\, 
        RDATA_IM0(42) => \RDATA_IM0[42]\, RDATA_IM0(41) => 
        \RDATA_IM0[41]\, RDATA_IM0(40) => \RDATA_IM0[40]\, 
        RDATA_IM0(39) => \RDATA_IM0[39]\, RDATA_IM0(38) => 
        \RDATA_IM0[38]\, RDATA_IM0(37) => \RDATA_IM0[37]\, 
        RDATA_IM0(36) => \RDATA_IM0[36]\, RDATA_IM0(35) => 
        \RDATA_IM0[35]\, RDATA_IM0(34) => \RDATA_IM0[34]\, 
        RDATA_IM0(33) => \RDATA_IM0[33]\, RDATA_IM0(32) => 
        \RDATA_IM0[32]\, RDATA_IM0(31) => \RDATA_IM0[31]\, 
        RDATA_IM0(30) => \RDATA_IM0[30]\, RDATA_IM0(29) => 
        \RDATA_IM0[29]\, RDATA_IM0(28) => \RDATA_IM0[28]\, 
        RDATA_IM0(27) => \RDATA_IM0[27]\, RDATA_IM0(26) => 
        \RDATA_IM0[26]\, RDATA_IM0(25) => \RDATA_IM0[25]\, 
        RDATA_IM0(24) => \RDATA_IM0[24]\, RDATA_IM0(23) => 
        \RDATA_IM0[23]\, RDATA_IM0(22) => \RDATA_IM0[22]\, 
        RDATA_IM0(21) => \RDATA_IM0[21]\, RDATA_IM0(20) => 
        \RDATA_IM0[20]\, RDATA_IM0(19) => \RDATA_IM0[19]\, 
        RDATA_IM0(18) => \RDATA_IM0[18]\, RDATA_IM0(17) => 
        \RDATA_IM0[17]\, RDATA_IM0(16) => \RDATA_IM0[16]\, 
        RDATA_IM0(15) => \RDATA_IM0[15]\, RDATA_IM0(14) => 
        \RDATA_IM0[14]\, RDATA_IM0(13) => \RDATA_IM0[13]\, 
        RDATA_IM0(12) => \RDATA_IM0[12]\, RDATA_IM0(11) => 
        \RDATA_IM0[11]\, RDATA_IM0(10) => \RDATA_IM0[10]\, 
        RDATA_IM0(9) => \RDATA_IM0[9]\, RDATA_IM0(8) => 
        \RDATA_IM0[8]\, RDATA_IM0(7) => \RDATA_IM0[7]\, 
        RDATA_IM0(6) => \RDATA_IM0[6]\, RDATA_IM0(5) => 
        \RDATA_IM0[5]\, RDATA_IM0(4) => \RDATA_IM0[4]\, 
        RDATA_IM0(3) => \RDATA_IM0[3]\, RDATA_IM0(2) => 
        \RDATA_IM0[2]\, RDATA_IM0(1) => \RDATA_IM0[1]\, 
        RDATA_IM0(0) => \RDATA_IM0[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1), 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1), AWADDR_MI0(27) => 
        \AWADDR_MI0[27]\, AWADDR_MI0(26) => \AWADDR_MI0[26]\, 
        AWADDR_MI0(25) => nc7, AWADDR_MI0(24) => nc6, 
        AWADDR_MI0(23) => \AWADDR_MI0[23]\, AWADDR_MI0(22) => 
        \AWADDR_MI0[22]\, AWADDR_MI0(21) => \AWADDR_MI0[21]\, 
        AWADDR_MI0(20) => \AWADDR_MI0[20]\, AWADDR_MI0(19) => 
        \AWADDR_MI0[19]\, AWADDR_MI0(18) => \AWADDR_MI0[18]\, 
        AWADDR_MI0(17) => \AWADDR_MI0[17]\, AWADDR_MI0(16) => 
        \AWADDR_MI0[16]\, AWADDR_MI0(15) => \AWADDR_MI0[15]\, 
        AWADDR_MI0(14) => \AWADDR_MI0[14]\, AWADDR_MI0(13) => 
        \AWADDR_MI0[13]\, AWADDR_MI0(12) => \AWADDR_MI0[12]\, 
        AWADDR_MI0(11) => \AWADDR_MI0[11]\, AWADDR_MI0(10) => 
        \AWADDR_MI0[10]\, AWADDR_MI0(9) => \AWADDR_MI0[9]\, 
        AWADDR_MI0(8) => \AWADDR_MI0[8]\, AWADDR_MI0(7) => 
        \AWADDR_MI0[7]\, AWADDR_MI0(6) => \AWADDR_MI0[6]\, 
        AWADDR_MI0(5) => \AWADDR_MI0[5]\, AWADDR_MI0(4) => 
        \AWADDR_MI0[4]\, AWADDR_MI0(3) => \AWADDR_MI0[3]\, 
        AWADDR_MI0(2) => \AWADDR_MI0[2]\, AWADDR_MI0(1) => 
        \AWADDR_MI0[1]\, ARADDR_MI0(27) => \ARADDR_MI0[27]\, 
        ARADDR_MI0(26) => \ARADDR_MI0[26]\, ARADDR_MI0(25) => 
        nc12, ARADDR_MI0(24) => nc5, ARADDR_MI0(23) => 
        \ARADDR_MI0[23]\, ARADDR_MI0(22) => \ARADDR_MI0[22]\, 
        ARADDR_MI0(21) => \ARADDR_MI0[21]\, ARADDR_MI0(20) => 
        \ARADDR_MI0[20]\, ARADDR_MI0(19) => \ARADDR_MI0[19]\, 
        ARADDR_MI0(18) => \ARADDR_MI0[18]\, ARADDR_MI0(17) => 
        \ARADDR_MI0[17]\, ARADDR_MI0(16) => \ARADDR_MI0[16]\, 
        ARADDR_MI0(15) => \ARADDR_MI0[15]\, ARADDR_MI0(14) => 
        \ARADDR_MI0[14]\, ARADDR_MI0(13) => \ARADDR_MI0[13]\, 
        ARADDR_MI0(12) => \ARADDR_MI0[12]\, ARADDR_MI0(11) => 
        \ARADDR_MI0[11]\, ARADDR_MI0(10) => \ARADDR_MI0[10]\, 
        ARADDR_MI0(9) => \ARADDR_MI0[9]\, ARADDR_MI0(8) => 
        \ARADDR_MI0[8]\, ARADDR_MI0(7) => \ARADDR_MI0[7]\, 
        ARADDR_MI0(6) => \ARADDR_MI0[6]\, ARADDR_MI0(5) => 
        \ARADDR_MI0[5]\, ARADDR_MI0(4) => \ARADDR_MI0[4]\, 
        ARADDR_MI0(3) => \ARADDR_MI0[3]\, ARADDR_MI0(2) => 
        \ARADDR_MI0[2]\, ARADDR_MI0(1) => \ARADDR_MI0[1]\, 
        ARSIZE_MI0(1) => \ARSIZE_MI0[1]\, ARSIZE_MI0(0) => 
        \ARSIZE_MI0[0]\, AWSIZE_MI0(1) => \AWSIZE_MI0[1]\, 
        AWSIZE_MI0(0) => \AWSIZE_MI0[0]\, WDATA_MI0(63) => 
        \WDATA_MI0[63]\, WDATA_MI0(62) => \WDATA_MI0[62]\, 
        WDATA_MI0(61) => \WDATA_MI0[61]\, WDATA_MI0(60) => 
        \WDATA_MI0[60]\, WDATA_MI0(59) => \WDATA_MI0[59]\, 
        WDATA_MI0(58) => \WDATA_MI0[58]\, WDATA_MI0(57) => 
        \WDATA_MI0[57]\, WDATA_MI0(56) => \WDATA_MI0[56]\, 
        WDATA_MI0(55) => \WDATA_MI0[55]\, WDATA_MI0(54) => 
        \WDATA_MI0[54]\, WDATA_MI0(53) => \WDATA_MI0[53]\, 
        WDATA_MI0(52) => \WDATA_MI0[52]\, WDATA_MI0(51) => 
        \WDATA_MI0[51]\, WDATA_MI0(50) => \WDATA_MI0[50]\, 
        WDATA_MI0(49) => \WDATA_MI0[49]\, WDATA_MI0(48) => 
        \WDATA_MI0[48]\, WDATA_MI0(47) => \WDATA_MI0[47]\, 
        WDATA_MI0(46) => \WDATA_MI0[46]\, WDATA_MI0(45) => 
        \WDATA_MI0[45]\, WDATA_MI0(44) => \WDATA_MI0[44]\, 
        WDATA_MI0(43) => \WDATA_MI0[43]\, WDATA_MI0(42) => 
        \WDATA_MI0[42]\, WDATA_MI0(41) => \WDATA_MI0[41]\, 
        WDATA_MI0(40) => \WDATA_MI0[40]\, WDATA_MI0(39) => 
        \WDATA_MI0[39]\, WDATA_MI0(38) => \WDATA_MI0[38]\, 
        WDATA_MI0(37) => \WDATA_MI0[37]\, WDATA_MI0(36) => 
        \WDATA_MI0[36]\, WDATA_MI0(35) => \WDATA_MI0[35]\, 
        WDATA_MI0(34) => \WDATA_MI0[34]\, WDATA_MI0(33) => 
        \WDATA_MI0[33]\, WDATA_MI0(32) => \WDATA_MI0[32]\, 
        WDATA_MI0(31) => \WDATA_MI0[31]\, WDATA_MI0(30) => 
        \WDATA_MI0[30]\, WDATA_MI0(29) => \WDATA_MI0[29]\, 
        WDATA_MI0(28) => \WDATA_MI0[28]\, WDATA_MI0(27) => 
        \WDATA_MI0[27]\, WDATA_MI0(26) => \WDATA_MI0[26]\, 
        WDATA_MI0(25) => \WDATA_MI0[25]\, WDATA_MI0(24) => 
        \WDATA_MI0[24]\, WDATA_MI0(23) => \WDATA_MI0[23]\, 
        WDATA_MI0(22) => \WDATA_MI0[22]\, WDATA_MI0(21) => 
        \WDATA_MI0[21]\, WDATA_MI0(20) => \WDATA_MI0[20]\, 
        WDATA_MI0(19) => \WDATA_MI0[19]\, WDATA_MI0(18) => 
        \WDATA_MI0[18]\, WDATA_MI0(17) => \WDATA_MI0[17]\, 
        WDATA_MI0(16) => \WDATA_MI0[16]\, WDATA_MI0(15) => 
        \WDATA_MI0[15]\, WDATA_MI0(14) => \WDATA_MI0[14]\, 
        WDATA_MI0(13) => \WDATA_MI0[13]\, WDATA_MI0(12) => 
        \WDATA_MI0[12]\, WDATA_MI0(11) => \WDATA_MI0[11]\, 
        WDATA_MI0(10) => \WDATA_MI0[10]\, WDATA_MI0(9) => 
        \WDATA_MI0[9]\, WDATA_MI0(8) => \WDATA_MI0[8]\, 
        WDATA_MI0(7) => \WDATA_MI0[7]\, WDATA_MI0(6) => 
        \WDATA_MI0[6]\, WDATA_MI0(5) => \WDATA_MI0[5]\, 
        WDATA_MI0(4) => \WDATA_MI0[4]\, WDATA_MI0(3) => 
        \WDATA_MI0[3]\, WDATA_MI0(2) => \WDATA_MI0[2]\, 
        WDATA_MI0(1) => \WDATA_MI0[1]\, WDATA_MI0(0) => 
        \WDATA_MI0[0]\, WSTRB_MI0(7) => \WSTRB_MI0[7]\, 
        WSTRB_MI0(6) => \WSTRB_MI0[6]\, WSTRB_MI0(5) => 
        \WSTRB_MI0[5]\, WSTRB_MI0(4) => \WSTRB_MI0[4]\, 
        WSTRB_MI0(3) => \WSTRB_MI0[3]\, WSTRB_MI0(2) => 
        \WSTRB_MI0[2]\, WSTRB_MI0(1) => \WSTRB_MI0[1]\, 
        WSTRB_MI0(0) => \WSTRB_MI0[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(63) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(63), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(31) => nc1, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(28) => nc9, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(21) => nc13, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(20) => nc8, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(19) => nc4, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0), axi_current_state_0
         => axi_current_state_0, axi_current_state_3 => 
        axi_current_state_3, ARBURST_MI0_0 => \ARBURST_MI0[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, AWLOCK_MI0_i_0 => 
        \AWLOCK_MI0_i[1]\, ARLOCK_MI0_i_0 => \ARLOCK_MI0_i[1]\, 
        ARREADY_IM0 => ARREADY_IM0, awaddr_awvalid_clr_d => 
        awaddr_awvalid_clr_d, RVALID_IM0 => RVALID_IM0, RLAST_IM0
         => RLAST_IM0, AWREADY_IM0 => AWREADY_IM0, WREADY_IM0 => 
        WREADY_IM0, COREAHBLTOAXI_0_AXIMasterIF_WVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, RREADY_MI0 => 
        RREADY_MI0, COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, araddr_arvalid_clr_d
         => araddr_arvalid_clr_d, BVALID_IM0 => BVALID_IM0, 
        m0_rd_end => m0_rd_end, 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, m0_wr_end => 
        m0_wr_end, COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\, 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, WVALID_MI0 => 
        WVALID_MI0, N_48 => N_48, AWVALID_MI0 => AWVALID_MI0, 
        ARVALID_MI0 => ARVALID_MI0, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, N_75_i => N_75_i, 
        N_135_i => N_135_i, N_136_i => N_136_i, N_137_i => 
        N_137_i, N_203_i => N_203_i, N_272_i => N_272_i, N_273_i
         => N_273_i, N_274_i => N_274_i, N_275_i => N_275_i, 
        N_276_i => N_276_i, N_277_i => N_277_i, N_382_i => 
        N_382_i, N_381_i => N_381_i, N_278_i => N_278_i, N_380_i
         => N_380_i, N_133_i => N_133_i, N_134_i => N_134_i, 
        N_195_i => N_195_i, N_197_i => N_197_i, N_200_i => 
        N_200_i, N_201_i => N_201_i, N_202_i => N_202_i, N_1452_i
         => N_1452_i, N_1451_i => N_1451_i, N_1450_i => N_1450_i, 
        N_1449_i => N_1449_i, N_1448_i => N_1448_i, N_1447_i => 
        N_1447_i, N_1446_i => N_1446_i, N_1445_i => N_1445_i, 
        wready_m_xhdl2 => wready_m_xhdl2, SDRCLK_c => SDRCLK_c, 
        MSS_READY => MSS_READY, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID);
    
    \L2.u_interconnect_ntom\ : axi_interconnect_ntom
      port map(AWSIZE_IS16_gated(1) => \AWSIZE_IS16_gated[1]\, 
        AWSIZE_IS16_gated(0) => \AWSIZE_IS16_gated[0]\, 
        AWADDR_MI0(27) => \AWADDR_MI0[27]\, AWADDR_MI0(26) => 
        \AWADDR_MI0[26]\, AWADDR_MI0(25) => nc11, AWADDR_MI0(24)
         => nc3, AWADDR_MI0(23) => \AWADDR_MI0[23]\, 
        AWADDR_MI0(22) => \AWADDR_MI0[22]\, AWADDR_MI0(21) => 
        \AWADDR_MI0[21]\, AWADDR_MI0(20) => \AWADDR_MI0[20]\, 
        AWADDR_MI0(19) => \AWADDR_MI0[19]\, AWADDR_MI0(18) => 
        \AWADDR_MI0[18]\, AWADDR_MI0(17) => \AWADDR_MI0[17]\, 
        AWADDR_MI0(16) => \AWADDR_MI0[16]\, AWADDR_MI0(15) => 
        \AWADDR_MI0[15]\, AWADDR_MI0(14) => \AWADDR_MI0[14]\, 
        AWADDR_MI0(13) => \AWADDR_MI0[13]\, AWADDR_MI0(12) => 
        \AWADDR_MI0[12]\, AWADDR_MI0(11) => \AWADDR_MI0[11]\, 
        AWADDR_MI0(10) => \AWADDR_MI0[10]\, AWADDR_MI0(9) => 
        \AWADDR_MI0[9]\, AWADDR_MI0(8) => \AWADDR_MI0[8]\, 
        AWADDR_MI0(7) => \AWADDR_MI0[7]\, AWADDR_MI0(6) => 
        \AWADDR_MI0[6]\, AWADDR_MI0(5) => \AWADDR_MI0[5]\, 
        AWADDR_MI0(4) => \AWADDR_MI0[4]\, AWADDR_MI0(3) => 
        \AWADDR_MI0[3]\, AWADDR_MI0(2) => \AWADDR_MI0[2]\, 
        AWADDR_MI0(1) => \AWADDR_MI0[1]\, AWADDR_IS16_gated(23)
         => \AWADDR_IS16_gated[23]\, AWADDR_IS16_gated(22) => 
        \AWADDR_IS16_gated[22]\, AWADDR_IS16_gated(21) => 
        \AWADDR_IS16_gated[21]\, AWADDR_IS16_gated(20) => 
        \AWADDR_IS16_gated[20]\, AWADDR_IS16_gated(19) => 
        \AWADDR_IS16_gated[19]\, AWADDR_IS16_gated(18) => 
        \AWADDR_IS16_gated[18]\, AWADDR_IS16_gated(17) => 
        \AWADDR_IS16_gated[17]\, AWADDR_IS16_gated(16) => 
        \AWADDR_IS16_gated[16]\, AWADDR_IS16_gated(15) => 
        \AWADDR_IS16_gated[15]\, AWADDR_IS16_gated(14) => 
        \AWADDR_IS16_gated[14]\, AWADDR_IS16_gated(13) => 
        \AWADDR_IS16_gated[13]\, AWADDR_IS16_gated(12) => 
        \AWADDR_IS16_gated[12]\, AWADDR_IS16_gated(11) => 
        \AWADDR_IS16_gated[11]\, AWADDR_IS16_gated(10) => 
        \AWADDR_IS16_gated[10]\, AWADDR_IS16_gated(9) => 
        \AWADDR_IS16_gated[9]\, AWADDR_IS16_gated(8) => 
        \AWADDR_IS16_gated[8]\, AWADDR_IS16_gated(7) => 
        \AWADDR_IS16_gated[7]\, AWADDR_IS16_gated(6) => 
        \AWADDR_IS16_gated[6]\, AWADDR_IS16_gated(5) => 
        \AWADDR_IS16_gated[5]\, AWADDR_IS16_gated(4) => 
        \AWADDR_IS16_gated[4]\, AWADDR_IS16_gated(3) => 
        \AWADDR_IS16_gated[3]\, AWADDR_IS16_gated(2) => 
        \AWADDR_IS16_gated[2]\, AWADDR_IS16_gated(1) => 
        \AWADDR_IS16_gated[1]\, AWSIZE_MI0(1) => \AWSIZE_MI0[1]\, 
        AWSIZE_MI0(0) => \AWSIZE_MI0[0]\, WDATA_MI0(63) => 
        \WDATA_MI0[63]\, WDATA_MI0(62) => \WDATA_MI0[62]\, 
        WDATA_MI0(61) => \WDATA_MI0[61]\, WDATA_MI0(60) => 
        \WDATA_MI0[60]\, WDATA_MI0(59) => \WDATA_MI0[59]\, 
        WDATA_MI0(58) => \WDATA_MI0[58]\, WDATA_MI0(57) => 
        \WDATA_MI0[57]\, WDATA_MI0(56) => \WDATA_MI0[56]\, 
        WDATA_MI0(55) => \WDATA_MI0[55]\, WDATA_MI0(54) => 
        \WDATA_MI0[54]\, WDATA_MI0(53) => \WDATA_MI0[53]\, 
        WDATA_MI0(52) => \WDATA_MI0[52]\, WDATA_MI0(51) => 
        \WDATA_MI0[51]\, WDATA_MI0(50) => \WDATA_MI0[50]\, 
        WDATA_MI0(49) => \WDATA_MI0[49]\, WDATA_MI0(48) => 
        \WDATA_MI0[48]\, WDATA_MI0(47) => \WDATA_MI0[47]\, 
        WDATA_MI0(46) => \WDATA_MI0[46]\, WDATA_MI0(45) => 
        \WDATA_MI0[45]\, WDATA_MI0(44) => \WDATA_MI0[44]\, 
        WDATA_MI0(43) => \WDATA_MI0[43]\, WDATA_MI0(42) => 
        \WDATA_MI0[42]\, WDATA_MI0(41) => \WDATA_MI0[41]\, 
        WDATA_MI0(40) => \WDATA_MI0[40]\, WDATA_MI0(39) => 
        \WDATA_MI0[39]\, WDATA_MI0(38) => \WDATA_MI0[38]\, 
        WDATA_MI0(37) => \WDATA_MI0[37]\, WDATA_MI0(36) => 
        \WDATA_MI0[36]\, WDATA_MI0(35) => \WDATA_MI0[35]\, 
        WDATA_MI0(34) => \WDATA_MI0[34]\, WDATA_MI0(33) => 
        \WDATA_MI0[33]\, WDATA_MI0(32) => \WDATA_MI0[32]\, 
        WDATA_MI0(31) => \WDATA_MI0[31]\, WDATA_MI0(30) => 
        \WDATA_MI0[30]\, WDATA_MI0(29) => \WDATA_MI0[29]\, 
        WDATA_MI0(28) => \WDATA_MI0[28]\, WDATA_MI0(27) => 
        \WDATA_MI0[27]\, WDATA_MI0(26) => \WDATA_MI0[26]\, 
        WDATA_MI0(25) => \WDATA_MI0[25]\, WDATA_MI0(24) => 
        \WDATA_MI0[24]\, WDATA_MI0(23) => \WDATA_MI0[23]\, 
        WDATA_MI0(22) => \WDATA_MI0[22]\, WDATA_MI0(21) => 
        \WDATA_MI0[21]\, WDATA_MI0(20) => \WDATA_MI0[20]\, 
        WDATA_MI0(19) => \WDATA_MI0[19]\, WDATA_MI0(18) => 
        \WDATA_MI0[18]\, WDATA_MI0(17) => \WDATA_MI0[17]\, 
        WDATA_MI0(16) => \WDATA_MI0[16]\, WDATA_MI0(15) => 
        \WDATA_MI0[15]\, WDATA_MI0(14) => \WDATA_MI0[14]\, 
        WDATA_MI0(13) => \WDATA_MI0[13]\, WDATA_MI0(12) => 
        \WDATA_MI0[12]\, WDATA_MI0(11) => \WDATA_MI0[11]\, 
        WDATA_MI0(10) => \WDATA_MI0[10]\, WDATA_MI0(9) => 
        \WDATA_MI0[9]\, WDATA_MI0(8) => \WDATA_MI0[8]\, 
        WDATA_MI0(7) => \WDATA_MI0[7]\, WDATA_MI0(6) => 
        \WDATA_MI0[6]\, WDATA_MI0(5) => \WDATA_MI0[5]\, 
        WDATA_MI0(4) => \WDATA_MI0[4]\, WDATA_MI0(3) => 
        \WDATA_MI0[3]\, WDATA_MI0(2) => \WDATA_MI0[2]\, 
        WDATA_MI0(1) => \WDATA_MI0[1]\, WDATA_MI0(0) => 
        \WDATA_MI0[0]\, WSTRB_MI0(7) => \WSTRB_MI0[7]\, 
        WSTRB_MI0(6) => \WSTRB_MI0[6]\, WSTRB_MI0(5) => 
        \WSTRB_MI0[5]\, WSTRB_MI0(4) => \WSTRB_MI0[4]\, 
        WSTRB_MI0(3) => \WSTRB_MI0[3]\, WSTRB_MI0(2) => 
        \WSTRB_MI0[2]\, WSTRB_MI0(1) => \WSTRB_MI0[1]\, 
        WSTRB_MI0(0) => \WSTRB_MI0[0]\, WDATA_IS16_gated(63) => 
        \WDATA_IS16_gated[63]\, WDATA_IS16_gated(62) => 
        \WDATA_IS16_gated[62]\, WDATA_IS16_gated(61) => 
        \WDATA_IS16_gated[61]\, WDATA_IS16_gated(60) => 
        \WDATA_IS16_gated[60]\, WDATA_IS16_gated(59) => 
        \WDATA_IS16_gated[59]\, WDATA_IS16_gated(58) => 
        \WDATA_IS16_gated[58]\, WDATA_IS16_gated(57) => 
        \WDATA_IS16_gated[57]\, WDATA_IS16_gated(56) => 
        \WDATA_IS16_gated[56]\, WDATA_IS16_gated(55) => 
        \WDATA_IS16_gated[55]\, WDATA_IS16_gated(54) => 
        \WDATA_IS16_gated[54]\, WDATA_IS16_gated(53) => 
        \WDATA_IS16_gated[53]\, WDATA_IS16_gated(52) => 
        \WDATA_IS16_gated[52]\, WDATA_IS16_gated(51) => 
        \WDATA_IS16_gated[51]\, WDATA_IS16_gated(50) => 
        \WDATA_IS16_gated[50]\, WDATA_IS16_gated(49) => 
        \WDATA_IS16_gated[49]\, WDATA_IS16_gated(48) => 
        \WDATA_IS16_gated[48]\, WDATA_IS16_gated(47) => 
        \WDATA_IS16_gated[47]\, WDATA_IS16_gated(46) => 
        \WDATA_IS16_gated[46]\, WDATA_IS16_gated(45) => 
        \WDATA_IS16_gated[45]\, WDATA_IS16_gated(44) => 
        \WDATA_IS16_gated[44]\, WDATA_IS16_gated(43) => 
        \WDATA_IS16_gated[43]\, WDATA_IS16_gated(42) => 
        \WDATA_IS16_gated[42]\, WDATA_IS16_gated(41) => 
        \WDATA_IS16_gated[41]\, WDATA_IS16_gated(40) => 
        \WDATA_IS16_gated[40]\, WDATA_IS16_gated(39) => 
        \WDATA_IS16_gated[39]\, WDATA_IS16_gated(38) => 
        \WDATA_IS16_gated[38]\, WDATA_IS16_gated(37) => 
        \WDATA_IS16_gated[37]\, WDATA_IS16_gated(36) => 
        \WDATA_IS16_gated[36]\, WDATA_IS16_gated(35) => 
        \WDATA_IS16_gated[35]\, WDATA_IS16_gated(34) => 
        \WDATA_IS16_gated[34]\, WDATA_IS16_gated(33) => 
        \WDATA_IS16_gated[33]\, WDATA_IS16_gated(32) => 
        \WDATA_IS16_gated[32]\, WDATA_IS16_gated(31) => 
        \WDATA_IS16_gated[31]\, WDATA_IS16_gated(30) => 
        \WDATA_IS16_gated[30]\, WDATA_IS16_gated(29) => 
        \WDATA_IS16_gated[29]\, WDATA_IS16_gated(28) => 
        \WDATA_IS16_gated[28]\, WDATA_IS16_gated(27) => 
        \WDATA_IS16_gated[27]\, WDATA_IS16_gated(26) => 
        \WDATA_IS16_gated[26]\, WDATA_IS16_gated(25) => 
        \WDATA_IS16_gated[25]\, WDATA_IS16_gated(24) => 
        \WDATA_IS16_gated[24]\, WDATA_IS16_gated(23) => 
        \WDATA_IS16_gated[23]\, WDATA_IS16_gated(22) => 
        \WDATA_IS16_gated[22]\, WDATA_IS16_gated(21) => 
        \WDATA_IS16_gated[21]\, WDATA_IS16_gated(20) => 
        \WDATA_IS16_gated[20]\, WDATA_IS16_gated(19) => 
        \WDATA_IS16_gated[19]\, WDATA_IS16_gated(18) => 
        \WDATA_IS16_gated[18]\, WDATA_IS16_gated(17) => 
        \WDATA_IS16_gated[17]\, WDATA_IS16_gated(16) => 
        \WDATA_IS16_gated[16]\, WDATA_IS16_gated(15) => 
        \WDATA_IS16_gated[15]\, WDATA_IS16_gated(14) => 
        \WDATA_IS16_gated[14]\, WDATA_IS16_gated(13) => 
        \WDATA_IS16_gated[13]\, WDATA_IS16_gated(12) => 
        \WDATA_IS16_gated[12]\, WDATA_IS16_gated(11) => 
        \WDATA_IS16_gated[11]\, WDATA_IS16_gated(10) => 
        \WDATA_IS16_gated[10]\, WDATA_IS16_gated(9) => 
        \WDATA_IS16_gated[9]\, WDATA_IS16_gated(8) => 
        \WDATA_IS16_gated[8]\, WDATA_IS16_gated(7) => 
        \WDATA_IS16_gated[7]\, WDATA_IS16_gated(6) => 
        \WDATA_IS16_gated[6]\, WDATA_IS16_gated(5) => 
        \WDATA_IS16_gated[5]\, WDATA_IS16_gated(4) => 
        \WDATA_IS16_gated[4]\, WDATA_IS16_gated(3) => 
        \WDATA_IS16_gated[3]\, WDATA_IS16_gated(2) => 
        \WDATA_IS16_gated[2]\, WDATA_IS16_gated(1) => 
        \WDATA_IS16_gated[1]\, WDATA_IS16_gated(0) => 
        \WDATA_IS16_gated[0]\, WSTRB_IS16_gated(7) => 
        \WSTRB_IS16_gated[7]\, WSTRB_IS16_gated(6) => 
        \WSTRB_IS16_gated[6]\, WSTRB_IS16_gated(5) => 
        \WSTRB_IS16_gated[5]\, WSTRB_IS16_gated(4) => 
        \WSTRB_IS16_gated[4]\, WSTRB_IS16_gated(3) => 
        \WSTRB_IS16_gated[3]\, WSTRB_IS16_gated(2) => 
        \WSTRB_IS16_gated[2]\, WSTRB_IS16_gated(1) => 
        \WSTRB_IS16_gated[1]\, WSTRB_IS16_gated(0) => 
        \WSTRB_IS16_gated[0]\, ARSIZE_IS16_gated(1) => 
        \ARSIZE_IS16_gated[1]\, ARSIZE_IS16_gated(0) => 
        \ARSIZE_IS16_gated[0]\, ARADDR_MI0(27) => 
        \ARADDR_MI0[27]\, ARADDR_MI0(26) => \ARADDR_MI0[26]\, 
        ARADDR_MI0(25) => nc10, ARADDR_MI0(24) => nc2, 
        ARADDR_MI0(23) => \ARADDR_MI0[23]\, ARADDR_MI0(22) => 
        \ARADDR_MI0[22]\, ARADDR_MI0(21) => \ARADDR_MI0[21]\, 
        ARADDR_MI0(20) => \ARADDR_MI0[20]\, ARADDR_MI0(19) => 
        \ARADDR_MI0[19]\, ARADDR_MI0(18) => \ARADDR_MI0[18]\, 
        ARADDR_MI0(17) => \ARADDR_MI0[17]\, ARADDR_MI0(16) => 
        \ARADDR_MI0[16]\, ARADDR_MI0(15) => \ARADDR_MI0[15]\, 
        ARADDR_MI0(14) => \ARADDR_MI0[14]\, ARADDR_MI0(13) => 
        \ARADDR_MI0[13]\, ARADDR_MI0(12) => \ARADDR_MI0[12]\, 
        ARADDR_MI0(11) => \ARADDR_MI0[11]\, ARADDR_MI0(10) => 
        \ARADDR_MI0[10]\, ARADDR_MI0(9) => \ARADDR_MI0[9]\, 
        ARADDR_MI0(8) => \ARADDR_MI0[8]\, ARADDR_MI0(7) => 
        \ARADDR_MI0[7]\, ARADDR_MI0(6) => \ARADDR_MI0[6]\, 
        ARADDR_MI0(5) => \ARADDR_MI0[5]\, ARADDR_MI0(4) => 
        \ARADDR_MI0[4]\, ARADDR_MI0(3) => \ARADDR_MI0[3]\, 
        ARADDR_MI0(2) => \ARADDR_MI0[2]\, ARADDR_MI0(1) => 
        \ARADDR_MI0[1]\, ARADDR_IS16_gated(23) => 
        \ARADDR_IS16_gated[23]\, ARADDR_IS16_gated(22) => 
        \ARADDR_IS16_gated[22]\, ARADDR_IS16_gated(21) => 
        \ARADDR_IS16_gated[21]\, ARADDR_IS16_gated(20) => 
        \ARADDR_IS16_gated[20]\, ARADDR_IS16_gated(19) => 
        \ARADDR_IS16_gated[19]\, ARADDR_IS16_gated(18) => 
        \ARADDR_IS16_gated[18]\, ARADDR_IS16_gated(17) => 
        \ARADDR_IS16_gated[17]\, ARADDR_IS16_gated(16) => 
        \ARADDR_IS16_gated[16]\, ARADDR_IS16_gated(15) => 
        \ARADDR_IS16_gated[15]\, ARADDR_IS16_gated(14) => 
        \ARADDR_IS16_gated[14]\, ARADDR_IS16_gated(13) => 
        \ARADDR_IS16_gated[13]\, ARADDR_IS16_gated(12) => 
        \ARADDR_IS16_gated[12]\, ARADDR_IS16_gated(11) => 
        \ARADDR_IS16_gated[11]\, ARADDR_IS16_gated(10) => 
        \ARADDR_IS16_gated[10]\, ARADDR_IS16_gated(9) => 
        \ARADDR_IS16_gated[9]\, ARADDR_IS16_gated(8) => 
        \ARADDR_IS16_gated[8]\, ARADDR_IS16_gated(7) => 
        \ARADDR_IS16_gated[7]\, ARADDR_IS16_gated(6) => 
        \ARADDR_IS16_gated[6]\, ARADDR_IS16_gated(5) => 
        \ARADDR_IS16_gated[5]\, ARADDR_IS16_gated(4) => 
        \ARADDR_IS16_gated[4]\, ARADDR_IS16_gated(3) => 
        \ARADDR_IS16_gated[3]\, ARADDR_IS16_gated(2) => 
        \ARADDR_IS16_gated[2]\, ARADDR_IS16_gated(1) => 
        \ARADDR_IS16_gated[1]\, ARSIZE_MI0(1) => \ARSIZE_MI0[1]\, 
        ARSIZE_MI0(0) => \ARSIZE_MI0[0]\, RDATA_IM0(63) => 
        \RDATA_IM0[63]\, RDATA_IM0(62) => \RDATA_IM0[62]\, 
        RDATA_IM0(61) => \RDATA_IM0[61]\, RDATA_IM0(60) => 
        \RDATA_IM0[60]\, RDATA_IM0(59) => \RDATA_IM0[59]\, 
        RDATA_IM0(58) => \RDATA_IM0[58]\, RDATA_IM0(57) => 
        \RDATA_IM0[57]\, RDATA_IM0(56) => \RDATA_IM0[56]\, 
        RDATA_IM0(55) => \RDATA_IM0[55]\, RDATA_IM0(54) => 
        \RDATA_IM0[54]\, RDATA_IM0(53) => \RDATA_IM0[53]\, 
        RDATA_IM0(52) => \RDATA_IM0[52]\, RDATA_IM0(51) => 
        \RDATA_IM0[51]\, RDATA_IM0(50) => \RDATA_IM0[50]\, 
        RDATA_IM0(49) => \RDATA_IM0[49]\, RDATA_IM0(48) => 
        \RDATA_IM0[48]\, RDATA_IM0(47) => \RDATA_IM0[47]\, 
        RDATA_IM0(46) => \RDATA_IM0[46]\, RDATA_IM0(45) => 
        \RDATA_IM0[45]\, RDATA_IM0(44) => \RDATA_IM0[44]\, 
        RDATA_IM0(43) => \RDATA_IM0[43]\, RDATA_IM0(42) => 
        \RDATA_IM0[42]\, RDATA_IM0(41) => \RDATA_IM0[41]\, 
        RDATA_IM0(40) => \RDATA_IM0[40]\, RDATA_IM0(39) => 
        \RDATA_IM0[39]\, RDATA_IM0(38) => \RDATA_IM0[38]\, 
        RDATA_IM0(37) => \RDATA_IM0[37]\, RDATA_IM0(36) => 
        \RDATA_IM0[36]\, RDATA_IM0(35) => \RDATA_IM0[35]\, 
        RDATA_IM0(34) => \RDATA_IM0[34]\, RDATA_IM0(33) => 
        \RDATA_IM0[33]\, RDATA_IM0(32) => \RDATA_IM0[32]\, 
        RDATA_IM0(31) => \RDATA_IM0[31]\, RDATA_IM0(30) => 
        \RDATA_IM0[30]\, RDATA_IM0(29) => \RDATA_IM0[29]\, 
        RDATA_IM0(28) => \RDATA_IM0[28]\, RDATA_IM0(27) => 
        \RDATA_IM0[27]\, RDATA_IM0(26) => \RDATA_IM0[26]\, 
        RDATA_IM0(25) => \RDATA_IM0[25]\, RDATA_IM0(24) => 
        \RDATA_IM0[24]\, RDATA_IM0(23) => \RDATA_IM0[23]\, 
        RDATA_IM0(22) => \RDATA_IM0[22]\, RDATA_IM0(21) => 
        \RDATA_IM0[21]\, RDATA_IM0(20) => \RDATA_IM0[20]\, 
        RDATA_IM0(19) => \RDATA_IM0[19]\, RDATA_IM0(18) => 
        \RDATA_IM0[18]\, RDATA_IM0(17) => \RDATA_IM0[17]\, 
        RDATA_IM0(16) => \RDATA_IM0[16]\, RDATA_IM0(15) => 
        \RDATA_IM0[15]\, RDATA_IM0(14) => \RDATA_IM0[14]\, 
        RDATA_IM0(13) => \RDATA_IM0[13]\, RDATA_IM0(12) => 
        \RDATA_IM0[12]\, RDATA_IM0(11) => \RDATA_IM0[11]\, 
        RDATA_IM0(10) => \RDATA_IM0[10]\, RDATA_IM0(9) => 
        \RDATA_IM0[9]\, RDATA_IM0(8) => \RDATA_IM0[8]\, 
        RDATA_IM0(7) => \RDATA_IM0[7]\, RDATA_IM0(6) => 
        \RDATA_IM0[6]\, RDATA_IM0(5) => \RDATA_IM0[5]\, 
        RDATA_IM0(4) => \RDATA_IM0[4]\, RDATA_IM0(3) => 
        \RDATA_IM0[3]\, RDATA_IM0(2) => \RDATA_IM0[2]\, 
        RDATA_IM0(1) => \RDATA_IM0[1]\, RDATA_IM0(0) => 
        \RDATA_IM0[0]\, COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, AWLOCK_MI0_i_0 => 
        \AWLOCK_MI0_i[1]\, ARBURST_IS16_gated_0 => 
        \ARBURST_IS16_gated[0]\, ARBURST_MI0_0 => 
        \ARBURST_MI0[0]\, ARLOCK_MI0_i_0 => \ARLOCK_MI0_i[1]\, 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        COREAXI_0_AXImslave16_RDATA_m_57, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        COREAXI_0_AXImslave16_RDATA_m_58, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        COREAXI_0_AXImslave16_RDATA_m_41, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        COREAXI_0_AXImslave16_RDATA_m_42, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        COREAXI_0_AXImslave16_RDATA_m_47, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        COREAXI_0_AXImslave16_RDATA_m_49, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        COREAXI_0_AXImslave16_RDATA_m_50, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        COREAXI_0_AXImslave16_RDATA_m_33, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        COREAXI_0_AXImslave16_RDATA_m_34, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        COREAXI_0_AXImslave16_RDATA_m_11, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        COREAXI_0_AXImslave16_RDATA_m_12, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        COREAXI_0_AXImslave16_RDATA_m_13, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        COREAXI_0_AXImslave16_RDATA_m_14, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        COREAXI_0_AXImslave16_RDATA_m_15, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        COREAXI_0_AXImslave16_RDATA_m_19, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        COREAXI_0_AXImslave16_RDATA_m_20, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        COREAXI_0_AXImslave16_RDATA_m_21, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        COREAXI_0_AXImslave16_RDATA_m_23, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        COREAXI_0_AXImslave16_RDATA_m_0, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        COREAXI_0_AXImslave16_RDATA_m_1, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        COREAXI_0_AXImslave16_RDATA_m_4, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        COREAXI_0_AXImslave16_RDATA_m_5, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        COREAXI_0_AXImslave16_RDATA_m_6, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        COREAXI_0_AXImslave16_RDATA_m_7, 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        COREAXI_0_AXImslave16_RDATA_m_8, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        COREAXI_0_AXImslave16_RDATA_m_9, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        COREAXI_0_AXImslave16_RDATA_m_10, 
        COREAXI_0_AXImslave16_RDATA_3 => 
        COREAXI_0_AXImslave16_RDATA_3, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        COREAXI_0_AXImslave16_RDATA_0, RDATA_reg_3 => RDATA_reg_3, 
        RDATA_reg_0 => RDATA_reg_0, axi_state_0 => axi_state_0, 
        AWREADY_IM0 => AWREADY_IM0, N_75_i => N_75_i, AWVALID_MI0
         => AWVALID_MI0, AWREADY_SI16 => AWREADY_SI16, m0_wr_end
         => m0_wr_end, WREADY_SI16 => WREADY_SI16, WVALID_MI0 => 
        WVALID_MI0, WREADY_IM0 => WREADY_IM0, ARREADY_IM0 => 
        ARREADY_IM0, COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, 
        COREAXI_0_AXImslave16_ARVALID => 
        \COREAXI_0_AXImslave16_ARVALID\, 
        COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, ARVALID_MI0 => ARVALID_MI0, 
        m0_rd_end => m0_rd_end, i22_mux_1_i => i22_mux_1_i, 
        i22_mux_0_i => i22_mux_0_i, i22_mux_i => i22_mux_i, 
        i17_mux_1_i => i17_mux_1_i, i17_mux_0_i => i17_mux_0_i, 
        i17_mux_i => i17_mux_i, N_3092_i => N_3092_i, N_3064_i
         => N_3064_i, i17_mux_2_i => i17_mux_2_i, N_8_i => N_8_i, 
        i22_mux_5_i => i22_mux_5_i, i22_mux_4_i => i22_mux_4_i, 
        i22_mux_3_i => i22_mux_3_i, i22_mux_2_i => i22_mux_2_i, 
        N_77_mux_i => N_77_mux_i, N_76_mux_i => N_76_mux_i, 
        N_75_mux_i => N_75_mux_i, N_69_mux_i => N_69_mux_i, 
        N_68_mux_i => N_68_mux_i, N_67_mux_i => N_67_mux_i, 
        N_3066_i => N_3066_i, N_3169_i => N_3169_i, N_3102_i => 
        N_3102_i, N_3100_i => N_3100_i, N_3098_i => N_3098_i, 
        N_3096_i => N_3096_i, N_3094_i => N_3094_i, N_72_mux_i
         => N_72_mux_i, N_71_mux_i => N_71_mux_i, N_70_mux_i => 
        N_70_mux_i, N_80_mux_i => N_80_mux_i, N_79_mux_i => 
        N_79_mux_i, N_78_mux_i => N_78_mux_i, N_39 => N_39, 
        N_3170_i => N_3170_i, RLAST_IM0 => RLAST_IM0, RVALID_IM0
         => RVALID_IM0, COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        \COREAHBLTOAXI_0_AXIMasterIF_RVALID\, N_23 => N_23, 
        N_3167_i => N_3167_i, N_74 => N_74, N_389 => N_389, 
        RREADY_MI0 => RREADY_MI0, N_3297 => N_3297, 
        COREAXI_0_AXImslave16_BVALID => 
        COREAXI_0_AXImslave16_BVALID, BVALID_IM0 => BVALID_IM0, 
        ARVALID_IS16 => ARVALID_IS16, AWVALID_IS16 => 
        AWVALID_IS16, WVALID_IS16 => WVALID_IS16, SDRCLK_c => 
        SDRCLK_c, MSS_READY => MSS_READY);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Synchronizer_AHBtoAXIHX is

    port( N_163_i            : in    std_logic;
          ahb_rd_req_sync    : out   std_logic;
          latch_ahb_sig      : in    std_logic;
          latch_ahb_sig_sync : out   std_logic;
          ahb_wr_done        : in    std_logic;
          wrch_fifo_wr_en_r  : out   std_logic;
          SDRCLK_c           : in    std_logic;
          ARESET_n           : in    std_logic;
          ahb_wr_done_sync   : out   std_logic
        );

end Synchronizer_AHBtoAXIHX;

architecture DEF_ARCH of Synchronizer_AHBtoAXIHX is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \wrch_fifo_wr_en_r\, GND_net_1, 
        \synchronizer_1[1]_net_1\, \synchronizer_3[1]_net_1\
         : std_logic;

begin 

    wrch_fifo_wr_en_r <= \wrch_fifo_wr_en_r\;

    \synchronizer_0[0]\ : SLE
      port map(D => \wrch_fifo_wr_en_r\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahb_wr_done_sync);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \synchronizer_3[1]\ : SLE
      port map(D => N_163_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_3[1]_net_1\);
    
    \synchronizer_3[0]\ : SLE
      port map(D => \synchronizer_3[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        ahb_rd_req_sync);
    
    \synchronizer_1[1]\ : SLE
      port map(D => latch_ahb_sig, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_1[1]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \synchronizer_1[0]\ : SLE
      port map(D => \synchronizer_1[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        latch_ahb_sig_sync);
    
    \synchronizer_0[1]\ : SLE
      port map(D => ahb_wr_done, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wrch_fifo_wr_en_r\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_wrch_ramHX is

    port( port_xhdl7        : out   std_logic_vector(63 downto 0);
          wrch_hwdata_r     : in    std_logic_vector(31 downto 0);
          wbinaddr          : in    std_logic_vector(3 downto 0);
          rbinaddr          : in    std_logic_vector(3 downto 0);
          wrch_fifo_wr_en_r : in    std_logic;
          fifo_full_xhdl2   : in    std_logic;
          wren_2            : in    std_logic;
          SDRCLK_c          : in    std_logic
        );

end CoreAHBLtoAXI_wrch_ramHX;

architecture DEF_ARCH of CoreAHBLtoAXI_wrch_ramHX is 

  component RAM64x18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_ADDR_CLK    : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ADDR_SRST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_ADDR_ARST_N : in    std_logic := 'U';
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_ADDR_EN     : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          B_ADDR_CLK    : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ADDR_SRST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_ADDR_ARST_N : in    std_logic := 'U';
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_ADDR_EN     : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_CLK         : in    std_logic := 'U';
          C_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          C_WEN         : in    std_logic := 'U';
          C_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_ADDR_LAT    : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_EN          : in    std_logic := 'U';
          B_ADDR_LAT    : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          C_EN          : in    std_logic := 'U';
          C_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1, mem2_mem2_0_0_we, 
        mem2_mem2_0_1_we, mem1_mem1_0_0_we, mem1_mem1_0_1_we
         : std_logic;
    signal nc47, nc34, nc70, nc60, nc74, nc64, nc9, nc13, nc23, 
        nc55, nc80, nc33, nc16, nc26, nc45, nc73, nc58, nc63, 
        nc27, nc17, nc36, nc48, nc37, nc5, nc52, nc76, nc51, nc66, 
        nc77, nc67, nc4, nc42, nc41, nc59, nc25, nc15, nc35, nc49, 
        nc28, nc18, nc75, nc65, nc38, nc1, nc2, nc50, nc22, nc12, 
        nc21, nc11, nc78, nc54, nc68, nc3, nc32, nc40, nc31, nc44, 
        nc7, nc72, nc6, nc71, nc62, nc61, nc19, nc29, nc53, nc39, 
        nc8, nc79, nc43, nc69, nc56, nc20, nc10, nc57, nc24, nc14, 
        nc46, nc30 : std_logic;

begin 


    mem2_mem2_0_1 : RAM64x18
      port map(A_DOUT(17) => nc47, A_DOUT(16) => nc34, A_DOUT(15)
         => port_xhdl7(63), A_DOUT(14) => port_xhdl7(62), 
        A_DOUT(13) => port_xhdl7(61), A_DOUT(12) => 
        port_xhdl7(60), A_DOUT(11) => port_xhdl7(59), A_DOUT(10)
         => port_xhdl7(58), A_DOUT(9) => port_xhdl7(57), 
        A_DOUT(8) => port_xhdl7(56), A_DOUT(7) => port_xhdl7(55), 
        A_DOUT(6) => port_xhdl7(54), A_DOUT(5) => port_xhdl7(53), 
        A_DOUT(4) => port_xhdl7(52), A_DOUT(3) => port_xhdl7(51), 
        A_DOUT(2) => port_xhdl7(50), A_DOUT(1) => port_xhdl7(49), 
        A_DOUT(0) => port_xhdl7(48), B_DOUT(17) => nc70, 
        B_DOUT(16) => nc60, B_DOUT(15) => nc74, B_DOUT(14) => 
        nc64, B_DOUT(13) => nc9, B_DOUT(12) => nc13, B_DOUT(11)
         => nc23, B_DOUT(10) => nc55, B_DOUT(9) => nc80, 
        B_DOUT(8) => nc33, B_DOUT(7) => nc16, B_DOUT(6) => nc26, 
        B_DOUT(5) => nc45, B_DOUT(4) => nc73, B_DOUT(3) => nc58, 
        B_DOUT(2) => nc63, B_DOUT(1) => nc27, B_DOUT(0) => nc17, 
        BUSY => OPEN, A_ADDR_CLK => SDRCLK_c, A_DOUT_CLK => 
        VCC_net_1, A_ADDR_SRST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_ADDR_ARST_N => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_ADDR_EN => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, A_ADDR(9)
         => GND_net_1, A_ADDR(8) => GND_net_1, A_ADDR(7) => 
        rbinaddr(3), A_ADDR(6) => rbinaddr(2), A_ADDR(5) => 
        rbinaddr(1), A_ADDR(4) => rbinaddr(0), A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, B_ADDR_CLK => SDRCLK_c, 
        B_DOUT_CLK => VCC_net_1, B_ADDR_SRST_N => VCC_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_ADDR_ARST_N => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_ADDR_EN => VCC_net_1, 
        B_DOUT_EN => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_ADDR(9) => GND_net_1, B_ADDR(8) => 
        GND_net_1, B_ADDR(7) => rbinaddr(3), B_ADDR(6) => 
        rbinaddr(2), B_ADDR(5) => rbinaddr(1), B_ADDR(4) => 
        rbinaddr(0), B_ADDR(3) => GND_net_1, B_ADDR(2) => 
        GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, 
        C_CLK => SDRCLK_c, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => wbinaddr(3), C_ADDR(6) => 
        wbinaddr(2), C_ADDR(5) => wbinaddr(1), C_ADDR(4) => 
        wbinaddr(0), C_ADDR(3) => GND_net_1, C_ADDR(2) => 
        GND_net_1, C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, 
        C_DIN(17) => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15)
         => wrch_hwdata_r(31), C_DIN(14) => wrch_hwdata_r(30), 
        C_DIN(13) => wrch_hwdata_r(29), C_DIN(12) => 
        wrch_hwdata_r(28), C_DIN(11) => wrch_hwdata_r(27), 
        C_DIN(10) => wrch_hwdata_r(26), C_DIN(9) => 
        wrch_hwdata_r(25), C_DIN(8) => wrch_hwdata_r(24), 
        C_DIN(7) => wrch_hwdata_r(23), C_DIN(6) => 
        wrch_hwdata_r(22), C_DIN(5) => wrch_hwdata_r(21), 
        C_DIN(4) => wrch_hwdata_r(20), C_DIN(3) => 
        wrch_hwdata_r(19), C_DIN(2) => wrch_hwdata_r(18), 
        C_DIN(1) => wrch_hwdata_r(17), C_DIN(0) => 
        wrch_hwdata_r(16), C_WEN => mem2_mem2_0_1_we, C_BLK(1)
         => VCC_net_1, C_BLK(0) => VCC_net_1, A_EN => VCC_net_1, 
        A_ADDR_LAT => GND_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => GND_net_1, 
        A_WIDTH(0) => GND_net_1, B_EN => GND_net_1, B_ADDR_LAT
         => GND_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        GND_net_1, C_EN => VCC_net_1, C_WIDTH(2) => VCC_net_1, 
        C_WIDTH(1) => GND_net_1, C_WIDTH(0) => GND_net_1, 
        SII_LOCK => GND_net_1);
    
    mem1_mem1_0_1_RNO : CFG3
      generic map(INIT => x"10")

      port map(A => fifo_full_xhdl2, B => wren_2, C => 
        wrch_fifo_wr_en_r, Y => mem1_mem1_0_1_we);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    mem2_mem2_0_0_RNO : CFG2
      generic map(INIT => x"2")

      port map(A => wren_2, B => fifo_full_xhdl2, Y => 
        mem2_mem2_0_0_we);
    
    mem1_mem1_0_1 : RAM64x18
      port map(A_DOUT(17) => nc36, A_DOUT(16) => nc48, A_DOUT(15)
         => port_xhdl7(31), A_DOUT(14) => port_xhdl7(30), 
        A_DOUT(13) => port_xhdl7(29), A_DOUT(12) => 
        port_xhdl7(28), A_DOUT(11) => port_xhdl7(27), A_DOUT(10)
         => port_xhdl7(26), A_DOUT(9) => port_xhdl7(25), 
        A_DOUT(8) => port_xhdl7(24), A_DOUT(7) => port_xhdl7(23), 
        A_DOUT(6) => port_xhdl7(22), A_DOUT(5) => port_xhdl7(21), 
        A_DOUT(4) => port_xhdl7(20), A_DOUT(3) => port_xhdl7(19), 
        A_DOUT(2) => port_xhdl7(18), A_DOUT(1) => port_xhdl7(17), 
        A_DOUT(0) => port_xhdl7(16), B_DOUT(17) => nc37, 
        B_DOUT(16) => nc5, B_DOUT(15) => nc52, B_DOUT(14) => nc76, 
        B_DOUT(13) => nc51, B_DOUT(12) => nc66, B_DOUT(11) => 
        nc77, B_DOUT(10) => nc67, B_DOUT(9) => nc4, B_DOUT(8) => 
        nc42, B_DOUT(7) => nc41, B_DOUT(6) => nc59, B_DOUT(5) => 
        nc25, B_DOUT(4) => nc15, B_DOUT(3) => nc35, B_DOUT(2) => 
        nc49, B_DOUT(1) => nc28, B_DOUT(0) => nc18, BUSY => OPEN, 
        A_ADDR_CLK => SDRCLK_c, A_DOUT_CLK => VCC_net_1, 
        A_ADDR_SRST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_ADDR_ARST_N => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, 
        A_ADDR_EN => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(1)
         => VCC_net_1, A_BLK(0) => VCC_net_1, A_ADDR(9) => 
        GND_net_1, A_ADDR(8) => GND_net_1, A_ADDR(7) => 
        rbinaddr(3), A_ADDR(6) => rbinaddr(2), A_ADDR(5) => 
        rbinaddr(1), A_ADDR(4) => rbinaddr(0), A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, B_ADDR_CLK => SDRCLK_c, 
        B_DOUT_CLK => VCC_net_1, B_ADDR_SRST_N => VCC_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_ADDR_ARST_N => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_ADDR_EN => VCC_net_1, 
        B_DOUT_EN => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_ADDR(9) => GND_net_1, B_ADDR(8) => 
        GND_net_1, B_ADDR(7) => rbinaddr(3), B_ADDR(6) => 
        rbinaddr(2), B_ADDR(5) => rbinaddr(1), B_ADDR(4) => 
        rbinaddr(0), B_ADDR(3) => GND_net_1, B_ADDR(2) => 
        GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, 
        C_CLK => SDRCLK_c, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => wbinaddr(3), C_ADDR(6) => 
        wbinaddr(2), C_ADDR(5) => wbinaddr(1), C_ADDR(4) => 
        wbinaddr(0), C_ADDR(3) => GND_net_1, C_ADDR(2) => 
        GND_net_1, C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, 
        C_DIN(17) => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15)
         => wrch_hwdata_r(31), C_DIN(14) => wrch_hwdata_r(30), 
        C_DIN(13) => wrch_hwdata_r(29), C_DIN(12) => 
        wrch_hwdata_r(28), C_DIN(11) => wrch_hwdata_r(27), 
        C_DIN(10) => wrch_hwdata_r(26), C_DIN(9) => 
        wrch_hwdata_r(25), C_DIN(8) => wrch_hwdata_r(24), 
        C_DIN(7) => wrch_hwdata_r(23), C_DIN(6) => 
        wrch_hwdata_r(22), C_DIN(5) => wrch_hwdata_r(21), 
        C_DIN(4) => wrch_hwdata_r(20), C_DIN(3) => 
        wrch_hwdata_r(19), C_DIN(2) => wrch_hwdata_r(18), 
        C_DIN(1) => wrch_hwdata_r(17), C_DIN(0) => 
        wrch_hwdata_r(16), C_WEN => mem1_mem1_0_1_we, C_BLK(1)
         => VCC_net_1, C_BLK(0) => VCC_net_1, A_EN => VCC_net_1, 
        A_ADDR_LAT => GND_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => GND_net_1, 
        A_WIDTH(0) => GND_net_1, B_EN => GND_net_1, B_ADDR_LAT
         => GND_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        VCC_net_1, B_WIDTH(1) => GND_net_1, B_WIDTH(0) => 
        GND_net_1, C_EN => VCC_net_1, C_WIDTH(2) => VCC_net_1, 
        C_WIDTH(1) => GND_net_1, C_WIDTH(0) => GND_net_1, 
        SII_LOCK => GND_net_1);
    
    mem2_mem2_0_1_RNO : CFG2
      generic map(INIT => x"2")

      port map(A => wren_2, B => fifo_full_xhdl2, Y => 
        mem2_mem2_0_1_we);
    
    mem2_mem2_0_0 : RAM64x18
      port map(A_DOUT(17) => nc75, A_DOUT(16) => nc65, A_DOUT(15)
         => port_xhdl7(47), A_DOUT(14) => port_xhdl7(46), 
        A_DOUT(13) => port_xhdl7(45), A_DOUT(12) => 
        port_xhdl7(44), A_DOUT(11) => port_xhdl7(43), A_DOUT(10)
         => port_xhdl7(42), A_DOUT(9) => port_xhdl7(41), 
        A_DOUT(8) => port_xhdl7(40), A_DOUT(7) => port_xhdl7(39), 
        A_DOUT(6) => port_xhdl7(38), A_DOUT(5) => port_xhdl7(37), 
        A_DOUT(4) => port_xhdl7(36), A_DOUT(3) => port_xhdl7(35), 
        A_DOUT(2) => port_xhdl7(34), A_DOUT(1) => port_xhdl7(33), 
        A_DOUT(0) => port_xhdl7(32), B_DOUT(17) => nc38, 
        B_DOUT(16) => nc1, B_DOUT(15) => nc2, B_DOUT(14) => nc50, 
        B_DOUT(13) => nc22, B_DOUT(12) => nc12, B_DOUT(11) => 
        nc21, B_DOUT(10) => nc11, B_DOUT(9) => nc78, B_DOUT(8)
         => nc54, B_DOUT(7) => nc68, B_DOUT(6) => nc3, B_DOUT(5)
         => nc32, B_DOUT(4) => nc40, B_DOUT(3) => nc31, B_DOUT(2)
         => nc44, B_DOUT(1) => nc7, B_DOUT(0) => nc72, BUSY => 
        OPEN, A_ADDR_CLK => SDRCLK_c, A_DOUT_CLK => VCC_net_1, 
        A_ADDR_SRST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_ADDR_ARST_N => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, 
        A_ADDR_EN => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(1)
         => VCC_net_1, A_BLK(0) => VCC_net_1, A_ADDR(9) => 
        GND_net_1, A_ADDR(8) => GND_net_1, A_ADDR(7) => 
        rbinaddr(3), A_ADDR(6) => rbinaddr(2), A_ADDR(5) => 
        rbinaddr(1), A_ADDR(4) => rbinaddr(0), A_ADDR(3) => 
        GND_net_1, A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, B_ADDR_CLK => SDRCLK_c, 
        B_DOUT_CLK => VCC_net_1, B_ADDR_SRST_N => VCC_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_ADDR_ARST_N => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_ADDR_EN => VCC_net_1, 
        B_DOUT_EN => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_ADDR(9) => GND_net_1, B_ADDR(8) => 
        GND_net_1, B_ADDR(7) => rbinaddr(3), B_ADDR(6) => 
        rbinaddr(2), B_ADDR(5) => rbinaddr(1), B_ADDR(4) => 
        rbinaddr(0), B_ADDR(3) => GND_net_1, B_ADDR(2) => 
        GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, 
        C_CLK => SDRCLK_c, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => wbinaddr(3), C_ADDR(6) => 
        wbinaddr(2), C_ADDR(5) => wbinaddr(1), C_ADDR(4) => 
        wbinaddr(0), C_ADDR(3) => GND_net_1, C_ADDR(2) => 
        GND_net_1, C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, 
        C_DIN(17) => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15)
         => wrch_hwdata_r(15), C_DIN(14) => wrch_hwdata_r(14), 
        C_DIN(13) => wrch_hwdata_r(13), C_DIN(12) => 
        wrch_hwdata_r(12), C_DIN(11) => wrch_hwdata_r(11), 
        C_DIN(10) => wrch_hwdata_r(10), C_DIN(9) => 
        wrch_hwdata_r(9), C_DIN(8) => wrch_hwdata_r(8), C_DIN(7)
         => wrch_hwdata_r(7), C_DIN(6) => wrch_hwdata_r(6), 
        C_DIN(5) => wrch_hwdata_r(5), C_DIN(4) => 
        wrch_hwdata_r(4), C_DIN(3) => wrch_hwdata_r(3), C_DIN(2)
         => wrch_hwdata_r(2), C_DIN(1) => wrch_hwdata_r(1), 
        C_DIN(0) => wrch_hwdata_r(0), C_WEN => mem2_mem2_0_0_we, 
        C_BLK(1) => VCC_net_1, C_BLK(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_ADDR_LAT => GND_net_1, A_DOUT_LAT => 
        VCC_net_1, A_WIDTH(2) => VCC_net_1, A_WIDTH(1) => 
        GND_net_1, A_WIDTH(0) => GND_net_1, B_EN => GND_net_1, 
        B_ADDR_LAT => GND_net_1, B_DOUT_LAT => VCC_net_1, 
        B_WIDTH(2) => VCC_net_1, B_WIDTH(1) => GND_net_1, 
        B_WIDTH(0) => GND_net_1, C_EN => VCC_net_1, C_WIDTH(2)
         => VCC_net_1, C_WIDTH(1) => GND_net_1, C_WIDTH(0) => 
        GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mem1_mem1_0_0_RNO : CFG3
      generic map(INIT => x"10")

      port map(A => fifo_full_xhdl2, B => wren_2, C => 
        wrch_fifo_wr_en_r, Y => mem1_mem1_0_0_we);
    
    mem1_mem1_0_0 : RAM64x18
      port map(A_DOUT(17) => nc6, A_DOUT(16) => nc71, A_DOUT(15)
         => port_xhdl7(15), A_DOUT(14) => port_xhdl7(14), 
        A_DOUT(13) => port_xhdl7(13), A_DOUT(12) => 
        port_xhdl7(12), A_DOUT(11) => port_xhdl7(11), A_DOUT(10)
         => port_xhdl7(10), A_DOUT(9) => port_xhdl7(9), A_DOUT(8)
         => port_xhdl7(8), A_DOUT(7) => port_xhdl7(7), A_DOUT(6)
         => port_xhdl7(6), A_DOUT(5) => port_xhdl7(5), A_DOUT(4)
         => port_xhdl7(4), A_DOUT(3) => port_xhdl7(3), A_DOUT(2)
         => port_xhdl7(2), A_DOUT(1) => port_xhdl7(1), A_DOUT(0)
         => port_xhdl7(0), B_DOUT(17) => nc62, B_DOUT(16) => nc61, 
        B_DOUT(15) => nc19, B_DOUT(14) => nc29, B_DOUT(13) => 
        nc53, B_DOUT(12) => nc39, B_DOUT(11) => nc8, B_DOUT(10)
         => nc79, B_DOUT(9) => nc43, B_DOUT(8) => nc69, B_DOUT(7)
         => nc56, B_DOUT(6) => nc20, B_DOUT(5) => nc10, B_DOUT(4)
         => nc57, B_DOUT(3) => nc24, B_DOUT(2) => nc14, B_DOUT(1)
         => nc46, B_DOUT(0) => nc30, BUSY => OPEN, A_ADDR_CLK => 
        SDRCLK_c, A_DOUT_CLK => VCC_net_1, A_ADDR_SRST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_ADDR_ARST_N => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_ADDR_EN => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(1) => VCC_net_1, 
        A_BLK(0) => VCC_net_1, A_ADDR(9) => GND_net_1, A_ADDR(8)
         => GND_net_1, A_ADDR(7) => rbinaddr(3), A_ADDR(6) => 
        rbinaddr(2), A_ADDR(5) => rbinaddr(1), A_ADDR(4) => 
        rbinaddr(0), A_ADDR(3) => GND_net_1, A_ADDR(2) => 
        GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, 
        B_ADDR_CLK => SDRCLK_c, B_DOUT_CLK => VCC_net_1, 
        B_ADDR_SRST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_ADDR_ARST_N => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, 
        B_ADDR_EN => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(1)
         => VCC_net_1, B_BLK(0) => VCC_net_1, B_ADDR(9) => 
        GND_net_1, B_ADDR(8) => GND_net_1, B_ADDR(7) => 
        rbinaddr(3), B_ADDR(6) => rbinaddr(2), B_ADDR(5) => 
        rbinaddr(1), B_ADDR(4) => rbinaddr(0), B_ADDR(3) => 
        GND_net_1, B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, C_CLK => SDRCLK_c, C_ADDR(9) => 
        GND_net_1, C_ADDR(8) => GND_net_1, C_ADDR(7) => 
        wbinaddr(3), C_ADDR(6) => wbinaddr(2), C_ADDR(5) => 
        wbinaddr(1), C_ADDR(4) => wbinaddr(0), C_ADDR(3) => 
        GND_net_1, C_ADDR(2) => GND_net_1, C_ADDR(1) => GND_net_1, 
        C_ADDR(0) => GND_net_1, C_DIN(17) => GND_net_1, C_DIN(16)
         => GND_net_1, C_DIN(15) => wrch_hwdata_r(15), C_DIN(14)
         => wrch_hwdata_r(14), C_DIN(13) => wrch_hwdata_r(13), 
        C_DIN(12) => wrch_hwdata_r(12), C_DIN(11) => 
        wrch_hwdata_r(11), C_DIN(10) => wrch_hwdata_r(10), 
        C_DIN(9) => wrch_hwdata_r(9), C_DIN(8) => 
        wrch_hwdata_r(8), C_DIN(7) => wrch_hwdata_r(7), C_DIN(6)
         => wrch_hwdata_r(6), C_DIN(5) => wrch_hwdata_r(5), 
        C_DIN(4) => wrch_hwdata_r(4), C_DIN(3) => 
        wrch_hwdata_r(3), C_DIN(2) => wrch_hwdata_r(2), C_DIN(1)
         => wrch_hwdata_r(1), C_DIN(0) => wrch_hwdata_r(0), C_WEN
         => mem1_mem1_0_0_we, C_BLK(1) => VCC_net_1, C_BLK(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_ADDR_LAT => GND_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => VCC_net_1, 
        A_WIDTH(1) => GND_net_1, A_WIDTH(0) => GND_net_1, B_EN
         => GND_net_1, B_ADDR_LAT => GND_net_1, B_DOUT_LAT => 
        VCC_net_1, B_WIDTH(2) => VCC_net_1, B_WIDTH(1) => 
        GND_net_1, B_WIDTH(0) => GND_net_1, C_EN => VCC_net_1, 
        C_WIDTH(2) => VCC_net_1, C_WIDTH(1) => GND_net_1, 
        C_WIDTH(0) => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_WRCHANNELFIFOHX is

    port( wrch_hwdata_r       : in    std_logic_vector(31 downto 0);
          masterAddrInProg_0  : in    std_logic;
          axi_current_state_0 : in    std_logic;
          valid_ahbcmd_i_o3_1 : in    std_logic;
          hsel2_0_a2_1        : in    std_logic;
          N_209               : out   std_logic;
          N_210               : out   std_logic;
          N_213               : out   std_logic;
          N_214               : out   std_logic;
          N_215               : out   std_logic;
          N_217               : out   std_logic;
          N_218               : out   std_logic;
          N_221               : out   std_logic;
          N_222               : out   std_logic;
          N_223               : out   std_logic;
          N_328               : out   std_logic;
          N_440               : out   std_logic;
          N_439               : out   std_logic;
          N_438               : out   std_logic;
          N_437               : out   std_logic;
          N_436               : out   std_logic;
          N_435               : out   std_logic;
          N_434               : out   std_logic;
          N_433               : out   std_logic;
          N_432               : out   std_logic;
          N_431               : out   std_logic;
          N_430               : out   std_logic;
          N_429               : out   std_logic;
          N_428               : out   std_logic;
          N_427               : out   std_logic;
          N_426               : out   std_logic;
          N_425               : out   std_logic;
          N_424               : out   std_logic;
          N_423               : out   std_logic;
          N_422               : out   std_logic;
          N_421               : out   std_logic;
          N_420               : out   std_logic;
          N_419               : out   std_logic;
          N_418               : out   std_logic;
          N_417               : out   std_logic;
          N_416               : out   std_logic;
          N_415               : out   std_logic;
          N_414               : out   std_logic;
          N_413               : out   std_logic;
          N_412               : out   std_logic;
          N_411               : out   std_logic;
          N_410               : out   std_logic;
          N_293               : out   std_logic;
          N_292               : out   std_logic;
          N_291               : out   std_logic;
          N_290               : out   std_logic;
          N_289               : out   std_logic;
          N_288               : out   std_logic;
          N_286               : out   std_logic;
          N_285               : out   std_logic;
          N_284               : out   std_logic;
          N_283               : out   std_logic;
          N_282               : out   std_logic;
          N_281               : out   std_logic;
          N_160               : out   std_logic;
          N_159               : out   std_logic;
          N_158               : out   std_logic;
          N_157               : out   std_logic;
          N_156               : out   std_logic;
          N_151               : out   std_logic;
          N_150               : out   std_logic;
          N_149               : out   std_logic;
          N_148               : out   std_logic;
          N_147               : out   std_logic;
          wrch_fifo_wr_en_r   : in    std_logic;
          ahb_busyidle_cyc    : in    std_logic;
          N_72_i              : in    std_logic;
          N_98                : in    std_logic;
          N_73_i_0            : in    std_logic;
          ahb_busyidle_cyc_i  : in    std_logic;
          SDRCLK_c            : in    std_logic;
          ARESET_n            : in    std_logic
        );

end CoreAHBLtoAXI_WRCHANNELFIFOHX;

architecture DEF_ARCH of CoreAHBLtoAXI_WRCHANNELFIFOHX is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CoreAHBLtoAXI_wrch_ramHX
    port( port_xhdl7        : out   std_logic_vector(63 downto 0);
          wrch_hwdata_r     : in    std_logic_vector(31 downto 0) := (others => 'U');
          wbinaddr          : in    std_logic_vector(3 downto 0) := (others => 'U');
          rbinaddr          : in    std_logic_vector(3 downto 0) := (others => 'U');
          wrch_fifo_wr_en_r : in    std_logic := 'U';
          fifo_full_xhdl2   : in    std_logic := 'U';
          wren_2            : in    std_logic := 'U';
          SDRCLK_c          : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal fifo_empty_xhdl3_0_N_2, fifo_empty_xhdl3_0_N_2_i, 
        \rsync2_wptr[32]_net_1\, VCC_net_1, 
        \rsync1_wptr[32]_net_1\, GND_net_1, 
        \rsync2_wptr[17]_net_1\, \rsync1_wptr[17]_net_1\, 
        \rsync2_wptr[18]_net_1\, \rsync1_wptr[18]_net_1\, 
        \rsync2_wptr[19]_net_1\, \rsync1_wptr[19]_net_1\, 
        \rsync2_wptr[20]_net_1\, \rsync1_wptr[20]_net_1\, 
        \rsync2_wptr[21]_net_1\, \rsync1_wptr[21]_net_1\, 
        \rsync2_wptr[22]_net_1\, \rsync1_wptr[22]_net_1\, 
        \rsync2_wptr[23]_net_1\, \rsync1_wptr[23]_net_1\, 
        \rsync2_wptr[24]_net_1\, \rsync1_wptr[24]_net_1\, 
        \rsync2_wptr[25]_net_1\, \rsync1_wptr[25]_net_1\, 
        \rsync2_wptr[26]_net_1\, \rsync1_wptr[26]_net_1\, 
        \rsync2_wptr[27]_net_1\, \rsync1_wptr[27]_net_1\, 
        \rsync2_wptr[28]_net_1\, \rsync1_wptr[28]_net_1\, 
        \rsync2_wptr[29]_net_1\, \rsync1_wptr[29]_net_1\, 
        \rsync2_wptr[30]_net_1\, \rsync1_wptr[30]_net_1\, 
        \rsync2_wptr[31]_net_1\, \rsync1_wptr[31]_net_1\, 
        \rsync2_wptr[2]_net_1\, \rsync1_wptr[2]_net_1\, 
        \rsync2_wptr[3]_net_1\, \rsync1_wptr[3]_net_1\, 
        \rsync2_wptr[4]_net_1\, \rsync1_wptr[4]_net_1\, 
        \rsync2_wptr[5]_net_1\, \rsync1_wptr[5]_net_1\, 
        \rsync2_wptr[6]_net_1\, \rsync1_wptr[6]_net_1\, 
        \rsync2_wptr[7]_net_1\, \rsync1_wptr[7]_net_1\, 
        \rsync2_wptr[8]_net_1\, \rsync1_wptr[8]_net_1\, 
        \rsync2_wptr[9]_net_1\, \rsync1_wptr[9]_net_1\, 
        \rsync2_wptr[10]_net_1\, \rsync1_wptr[10]_net_1\, 
        \rsync2_wptr[11]_net_1\, \rsync1_wptr[11]_net_1\, 
        \rsync2_wptr[12]_net_1\, \rsync1_wptr[12]_net_1\, 
        \rsync2_wptr[13]_net_1\, \rsync1_wptr[13]_net_1\, 
        \rsync2_wptr[14]_net_1\, \rsync1_wptr[14]_net_1\, 
        \rsync2_wptr[15]_net_1\, \rsync1_wptr[15]_net_1\, 
        \rsync2_wptr[16]_net_1\, \rsync1_wptr[16]_net_1\, 
        \wsync2_rptr[20]_net_1\, \wsync1_rptr[20]_net_1\, 
        \wsync2_rptr[21]_net_1\, \wsync1_rptr[21]_net_1\, 
        \wsync2_rptr[22]_net_1\, \wsync1_rptr[22]_net_1\, 
        \wsync2_rptr[23]_net_1\, \wsync1_rptr[23]_net_1\, 
        \wsync2_rptr[24]_net_1\, \wsync1_rptr[24]_net_1\, 
        \wsync2_rptr[25]_net_1\, \wsync1_rptr[25]_net_1\, 
        \wsync2_rptr[26]_net_1\, \wsync1_rptr[26]_net_1\, 
        \wsync2_rptr[27]_net_1\, \wsync1_rptr[27]_net_1\, 
        \wsync2_rptr[28]_net_1\, \wsync1_rptr[28]_net_1\, 
        \wsync2_rptr[29]_net_1\, \wsync1_rptr[29]_net_1\, 
        \wsync2_rptr[30]_net_1\, \wsync1_rptr[30]_net_1\, 
        \wsync2_rptr[31]_net_1\, \wsync1_rptr[31]_net_1\, 
        \wsync2_rptr[32]_net_1\, \wsync1_rptr[32]_net_1\, 
        \rsync2_wptr[0]_net_1\, \rsync1_wptr[0]_net_1\, 
        \rsync2_wptr[1]_net_1\, \rsync1_wptr[1]_net_1\, 
        \wsync2_rptr[5]_net_1\, \wsync1_rptr[5]_net_1\, 
        \wsync2_rptr[6]_net_1\, \wsync1_rptr[6]_net_1\, 
        \wsync2_rptr[7]_net_1\, \wsync1_rptr[7]_net_1\, 
        \wsync2_rptr[8]_net_1\, \wsync1_rptr[8]_net_1\, 
        \wsync2_rptr[9]_net_1\, \wsync1_rptr[9]_net_1\, 
        \wsync2_rptr[10]_net_1\, \wsync1_rptr[10]_net_1\, 
        \wsync2_rptr[11]_net_1\, \wsync1_rptr[11]_net_1\, 
        \wsync2_rptr[12]_net_1\, \wsync1_rptr[12]_net_1\, 
        \wsync2_rptr[13]_net_1\, \wsync1_rptr[13]_net_1\, 
        \wsync2_rptr[14]_net_1\, \wsync1_rptr[14]_net_1\, 
        \wsync2_rptr[15]_net_1\, \wsync1_rptr[15]_net_1\, 
        \wsync2_rptr[16]_net_1\, \wsync1_rptr[16]_net_1\, 
        \wsync2_rptr[17]_net_1\, \wsync1_rptr[17]_net_1\, 
        \wsync2_rptr[18]_net_1\, \wsync1_rptr[18]_net_1\, 
        \wsync2_rptr[19]_net_1\, \wsync1_rptr[19]_net_1\, 
        \waddr_gray[23]_net_1\, \waddr_gray[24]_net_1\, 
        \waddr_gray[25]_net_1\, \waddr_gray[26]_net_1\, 
        \waddr_gray[27]_net_1\, \waddr_gray[28]_net_1\, 
        \waddr_gray[29]_net_1\, \waddr_gray[30]_net_1\, 
        \waddr_gray[31]_net_1\, \waddr_gray[32]_net_1\, 
        \wsync2_rptr[0]_net_1\, \wsync1_rptr[0]_net_1\, 
        \wsync2_rptr[1]_net_1\, \wsync1_rptr[1]_net_1\, 
        \wsync2_rptr[2]_net_1\, \wsync1_rptr[2]_net_1\, 
        \wsync2_rptr[3]_net_1\, \wsync1_rptr[3]_net_1\, 
        \wsync2_rptr[4]_net_1\, \wsync1_rptr[4]_net_1\, 
        \waddr_gray[8]_net_1\, \waddr_gray[9]_net_1\, 
        \waddr_gray[10]_net_1\, \waddr_gray[11]_net_1\, 
        \waddr_gray[12]_net_1\, \waddr_gray[13]_net_1\, 
        \waddr_gray[14]_net_1\, \waddr_gray[15]_net_1\, 
        \waddr_gray[16]_net_1\, \waddr_gray[17]_net_1\, 
        \waddr_gray[18]_net_1\, \waddr_gray[19]_net_1\, 
        \waddr_gray[20]_net_1\, \waddr_gray[21]_net_1\, 
        \waddr_gray[22]_net_1\, \raddr_gray[26]_net_1\, 
        \raddr_gray[27]_net_1\, \raddr_gray[28]_net_1\, 
        \raddr_gray[29]_net_1\, \raddr_gray[30]_net_1\, 
        \raddr_gray[31]_net_1\, \raddr_gray[32]_net_1\, 
        \waddr_gray[0]_net_1\, \waddr_gray[1]_net_1\, 
        \waddr_gray[2]_net_1\, \waddr_gray[3]_net_1\, 
        \waddr_gray[4]_net_1\, \waddr_gray[5]_net_1\, 
        \waddr_gray[6]_net_1\, \waddr_gray[7]_net_1\, 
        \raddr_gray[11]_net_1\, \raddr_gray[12]_net_1\, 
        \raddr_gray[13]_net_1\, \raddr_gray[14]_net_1\, 
        \raddr_gray[15]_net_1\, \raddr_gray[16]_net_1\, 
        \raddr_gray[17]_net_1\, \raddr_gray[18]_net_1\, 
        \raddr_gray[19]_net_1\, \raddr_gray[20]_net_1\, 
        \raddr_gray[21]_net_1\, \raddr_gray[22]_net_1\, 
        \raddr_gray[23]_net_1\, \raddr_gray[24]_net_1\, 
        \raddr_gray[25]_net_1\, \wgraynext[29]_net_1\, 
        \wgraynext[30]_net_1\, \wgraynext[31]_net_1\, 
        \wbinaddr_RNIKGF6A_S[32]\, \raddr_gray[0]_net_1\, 
        \raddr_gray[1]_net_1\, \raddr_gray[2]_net_1\, 
        \raddr_gray[3]_net_1\, \raddr_gray[4]_net_1\, 
        \raddr_gray[5]_net_1\, \raddr_gray[6]_net_1\, 
        \raddr_gray[7]_net_1\, \raddr_gray[8]_net_1\, 
        \raddr_gray[9]_net_1\, \raddr_gray[10]_net_1\, 
        \wgraynext[14]_net_1\, \wgraynext[15]_net_1\, 
        \wgraynext[16]_net_1\, \wgraynext[17]_net_1\, 
        \wgraynext[18]_net_1\, \wgraynext[19]_net_1\, 
        \wgraynext[20]_net_1\, \wgraynext[21]_net_1\, 
        \wgraynext[22]_net_1\, \wgraynext[23]_net_1\, 
        \wgraynext[24]_net_1\, \wgraynext[25]_net_1\, 
        \wgraynext[26]_net_1\, \wgraynext[27]_net_1\, 
        \wgraynext[28]_net_1\, \wbinaddr[32]_net_1\, 
        \wbinaddr_2[32]\, \wgraynext[0]_net_1\, 
        \wgraynext[1]_net_1\, \wgraynext[2]_net_1\, 
        \wgraynext[3]_net_1\, \wgraynext[4]_net_1\, 
        \wgraynext[5]_net_1\, \wgraynext[6]_net_1\, 
        \wgraynext[7]_net_1\, \wgraynext[8]_net_1\, 
        \wgraynext[9]_net_1\, \wgraynext[10]_net_1\, 
        \wgraynext[11]_net_1\, \wgraynext[12]_net_1\, 
        \wgraynext[13]_net_1\, \wbinaddr[17]_net_1\, 
        \wbinaddr_2[17]\, \wbinaddr[18]_net_1\, \wbinaddr_2[18]\, 
        \wbinaddr[19]_net_1\, \wbinaddr_2[19]\, 
        \wbinaddr[20]_net_1\, \wbinaddr_2[20]\, 
        \wbinaddr[21]_net_1\, \wbinaddr_2[21]\, 
        \wbinaddr[22]_net_1\, \wbinaddr_2[22]\, 
        \wbinaddr[23]_net_1\, \wbinaddr_2[23]\, 
        \wbinaddr[24]_net_1\, \wbinaddr_2[24]\, 
        \wbinaddr[25]_net_1\, \wbinaddr_2[25]\, 
        \wbinaddr[26]_net_1\, \wbinaddr_2[26]\, 
        \wbinaddr[27]_net_1\, \wbinaddr_2[27]\, 
        \wbinaddr[28]_net_1\, \wbinaddr_2[28]\, 
        \wbinaddr[29]_net_1\, \wbinaddr_2[29]\, 
        \wbinaddr[30]_net_1\, \wbinaddr_2[30]\, 
        \wbinaddr[31]_net_1\, \wbinaddr_2[31]\, 
        \wbinaddr[2]_net_1\, \wbinaddr_2[2]\, \wbinaddr[3]_net_1\, 
        \wbinaddr_2[3]\, \wbinaddr[4]_net_1\, \wbinaddr_2[4]\, 
        \wbinaddr[5]_net_1\, \wbinaddr_2[5]\, \wbinaddr[6]_net_1\, 
        \wbinaddr_2[6]\, \wbinaddr[7]_net_1\, \wbinaddr_2[7]\, 
        \wbinaddr[8]_net_1\, \wbinaddr_2[8]\, \wbinaddr[9]_net_1\, 
        \wbinaddr_2[9]\, \wbinaddr[10]_net_1\, \wbinaddr_2[10]\, 
        \wbinaddr[11]_net_1\, \wbinaddr_2[11]\, 
        \wbinaddr[12]_net_1\, \wbinaddr_2[12]\, 
        \wbinaddr[13]_net_1\, \wbinaddr_2[13]\, 
        \wbinaddr[14]_net_1\, \wbinaddr_2[14]\, 
        \wbinaddr[15]_net_1\, \wbinaddr_2[15]\, 
        \wbinaddr[16]_net_1\, \wbinaddr_2[16]\, 
        \rgraynext[20]_net_1\, \rgraynext[21]_net_1\, 
        \rgraynext[22]_net_1\, \rgraynext[23]_net_1\, 
        \rgraynext[24]_net_1\, \rgraynext[25]_net_1\, 
        \rgraynext[26]_net_1\, \rgraynext[27]_net_1\, 
        \rgraynext[28]_net_1\, \rgraynext[29]_net_1\, 
        \rgraynext[30]_net_1\, \rgraynext[31]_net_1\, 
        \rbinaddr_RNI79FFG_S[32]\, \wbinaddr[0]_net_1\, 
        \wbinaddr_2[0]\, \wbinaddr[1]_net_1\, \wbinaddr_2[1]\, 
        \rgraynext[5]_net_1\, \rgraynext[6]_net_1\, 
        \rgraynext[7]_net_1\, \rgraynext[8]_net_1\, 
        \rgraynext[9]_net_1\, \rgraynext[10]_net_1\, 
        \rgraynext[11]_net_1\, \rgraynext[12]_net_1\, 
        \rgraynext[13]_net_1\, \rgraynext[14]_net_1\, 
        \rgraynext[15]_net_1\, \rgraynext[16]_net_1\, 
        \rgraynext[17]_net_1\, \rgraynext[18]_net_1\, 
        \rgraynext[19]_net_1\, \rbinaddr[23]_net_1\, 
        \rbinaddr_3[23]\, \rbinaddr[24]_net_1\, \rbinaddr_3[24]\, 
        \rbinaddr[25]_net_1\, \rbinaddr_3[25]\, 
        \rbinaddr[26]_net_1\, \rbinaddr_3[26]\, 
        \rbinaddr[27]_net_1\, \rbinaddr_3[27]\, 
        \rbinaddr[28]_net_1\, \rbinaddr_3[28]\, 
        \rbinaddr[29]_net_1\, \rbinaddr_3[29]\, 
        \rbinaddr[30]_net_1\, \rbinaddr_3[30]\, 
        \rbinaddr[31]_net_1\, \rbinaddr_3[31]\, 
        \rbinaddr[32]_net_1\, \rbinaddr_3[32]\, 
        \rgraynext[0]_net_1\, \rgraynext[1]_net_1\, 
        \rgraynext[2]_net_1\, \rgraynext[3]_net_1\, 
        \rgraynext[4]_net_1\, \rbinaddr[8]_net_1\, 
        \rbinaddr_3[8]\, \rbinaddr[9]_net_1\, \rbinaddr_3[9]\, 
        \rbinaddr[10]_net_1\, \rbinaddr_3[10]\, 
        \rbinaddr[11]_net_1\, \rbinaddr_3[11]\, 
        \rbinaddr[12]_net_1\, \rbinaddr_3[12]\, 
        \rbinaddr[13]_net_1\, \rbinaddr_3[13]\, 
        \rbinaddr[14]_net_1\, \rbinaddr_3[14]\, 
        \rbinaddr[15]_net_1\, \rbinaddr_3[15]\, 
        \rbinaddr[16]_net_1\, \rbinaddr_3[16]\, 
        \rbinaddr[17]_net_1\, \rbinaddr_3[17]\, 
        \rbinaddr[18]_net_1\, \rbinaddr_3[18]\, 
        \rbinaddr[19]_net_1\, \rbinaddr_3[19]\, 
        \rbinaddr[20]_net_1\, \rbinaddr_3[20]\, 
        \rbinaddr[21]_net_1\, \rbinaddr_3[21]\, 
        \rbinaddr[22]_net_1\, \rbinaddr_3[22]\, 
        \rddata_r[57]_net_1\, \port_xhdl7[57]\, \rdinr_d\, 
        \rddata_r[58]_net_1\, \port_xhdl7[58]\, 
        \rddata_r[59]_net_1\, \port_xhdl7[59]\, 
        \rddata_r[60]_net_1\, \port_xhdl7[60]\, 
        \rddata_r[61]_net_1\, \port_xhdl7[61]\, 
        \rddata_r[62]_net_1\, \port_xhdl7[62]\, 
        \rddata_r[63]_net_1\, \port_xhdl7[63]\, 
        \rbinaddr[0]_net_1\, \rbinaddr_3[0]\, \rbinaddr[1]_net_1\, 
        \rbinaddr_3[1]\, \rbinaddr[2]_net_1\, \rbinaddr_3[2]\, 
        \rbinaddr[3]_net_1\, \rbinaddr_3[3]\, \rbinaddr[4]_net_1\, 
        \rbinaddr_3[4]\, \rbinaddr[5]_net_1\, \rbinaddr_3[5]\, 
        \rbinaddr[6]_net_1\, \rbinaddr_3[6]\, \rbinaddr[7]_net_1\, 
        \rbinaddr_3[7]\, \rddata_r[42]_net_1\, \port_xhdl7[42]\, 
        \rddata_r[43]_net_1\, \port_xhdl7[43]\, 
        \rddata_r[44]_net_1\, \port_xhdl7[44]\, 
        \rddata_r[45]_net_1\, \port_xhdl7[45]\, 
        \rddata_r[46]_net_1\, \port_xhdl7[46]\, 
        \rddata_r[47]_net_1\, \port_xhdl7[47]\, 
        \rddata_r[48]_net_1\, \port_xhdl7[48]\, 
        \rddata_r[49]_net_1\, \port_xhdl7[49]\, 
        \rddata_r[50]_net_1\, \port_xhdl7[50]\, 
        \rddata_r[51]_net_1\, \port_xhdl7[51]\, 
        \rddata_r[52]_net_1\, \port_xhdl7[52]\, 
        \rddata_r[53]_net_1\, \port_xhdl7[53]\, 
        \rddata_r[54]_net_1\, \port_xhdl7[54]\, 
        \rddata_r[55]_net_1\, \port_xhdl7[55]\, 
        \rddata_r[56]_net_1\, \port_xhdl7[56]\, 
        \rddata_r[27]_net_1\, \port_xhdl7[27]\, 
        \rddata_r[28]_net_1\, \port_xhdl7[28]\, 
        \rddata_r[29]_net_1\, \port_xhdl7[29]\, 
        \rddata_r[30]_net_1\, \port_xhdl7[30]\, 
        \rddata_r[31]_net_1\, \port_xhdl7[31]\, 
        \rddata_r[32]_net_1\, \port_xhdl7[32]\, 
        \rddata_r[33]_net_1\, \port_xhdl7[33]\, 
        \rddata_r[34]_net_1\, \port_xhdl7[34]\, 
        \rddata_r[35]_net_1\, \port_xhdl7[35]\, 
        \rddata_r[36]_net_1\, \port_xhdl7[36]\, 
        \rddata_r[37]_net_1\, \port_xhdl7[37]\, 
        \rddata_r[38]_net_1\, \port_xhdl7[38]\, 
        \rddata_r[39]_net_1\, \port_xhdl7[39]\, 
        \rddata_r[40]_net_1\, \port_xhdl7[40]\, 
        \rddata_r[41]_net_1\, \port_xhdl7[41]\, 
        \rddata_r[12]_net_1\, \port_xhdl7[12]\, 
        \rddata_r[13]_net_1\, \port_xhdl7[13]\, 
        \rddata_r[14]_net_1\, \port_xhdl7[14]\, 
        \rddata_r[15]_net_1\, \port_xhdl7[15]\, 
        \rddata_r[16]_net_1\, \port_xhdl7[16]\, 
        \rddata_r[17]_net_1\, \port_xhdl7[17]\, 
        \rddata_r[18]_net_1\, \port_xhdl7[18]\, 
        \rddata_r[19]_net_1\, \port_xhdl7[19]\, 
        \rddata_r[20]_net_1\, \port_xhdl7[20]\, 
        \rddata_r[21]_net_1\, \port_xhdl7[21]\, 
        \rddata_r[22]_net_1\, \port_xhdl7[22]\, 
        \rddata_r[23]_net_1\, \port_xhdl7[23]\, 
        \rddata_r[24]_net_1\, \port_xhdl7[24]\, 
        \rddata_r[25]_net_1\, \port_xhdl7[25]\, 
        \rddata_r[26]_net_1\, \port_xhdl7[26]\, 
        \rddata_r[0]_net_1\, \port_xhdl7[0]\, \rddata_r[1]_net_1\, 
        \port_xhdl7[1]\, \rddata_r[2]_net_1\, \port_xhdl7[2]\, 
        \rddata_r[3]_net_1\, \port_xhdl7[3]\, \rddata_r[4]_net_1\, 
        \port_xhdl7[4]\, \rddata_r[5]_net_1\, \port_xhdl7[5]\, 
        \rddata_r[6]_net_1\, \port_xhdl7[6]\, \rddata_r[7]_net_1\, 
        \port_xhdl7[7]\, \rddata_r[8]_net_1\, \port_xhdl7[8]\, 
        \rddata_r[9]_net_1\, \port_xhdl7[9]\, 
        \rddata_r[10]_net_1\, \port_xhdl7[10]\, 
        \rddata_r[11]_net_1\, \port_xhdl7[11]\, \wren_2\, 
        \wren_1\, \fifo_empty_xhdl3\, \fifo_full_xhdl2\, 
        \un9_writefull\, un3_rbinnext_cry_0_cy, 
        un3_rbinnext_cry_0, \rbinaddr_RNI6KBL1_S[0]\, 
        un3_rbinnext_cry_1, \rbinaddr_RNI32A52_S[1]\, 
        un3_rbinnext_cry_2, \rbinaddr_RNI1H8L2_S[2]\, 
        un3_rbinnext_cry_3, \rbinaddr_RNI01753_S[3]\, 
        un3_rbinnext_cry_4, \rbinaddr_RNI0I5L3_S[4]\, 
        un3_rbinnext_cry_5, \rbinaddr_RNI14454_S[5]\, 
        un3_rbinnext_cry_6, \rbinaddr_RNI3N2L4_S[6]\, 
        un3_rbinnext_cry_7, \rbinaddr_RNI6B155_S[7]\, 
        un3_rbinnext_cry_8, \rbinaddr_RNIA00L5_S[8]\, 
        un3_rbinnext_cry_9, \rbinaddr_RNIFMU46_S[9]\, 
        un3_rbinnext_cry_10, \rbinaddr_RNISL9J6_S[10]\, 
        un3_rbinnext_cry_11, \rbinaddr_RNIAMK17_S[11]\, 
        un3_rbinnext_cry_12, \rbinaddr_RNIPNVF7_S[12]\, 
        un3_rbinnext_cry_13, \rbinaddr_RNI9QAU7_S[13]\, 
        un3_rbinnext_cry_14, \rbinaddr_RNIQTLC8_S[14]\, 
        un3_rbinnext_cry_15, \rbinaddr_RNIC21R8_S[15]\, 
        un3_rbinnext_cry_16, \rbinaddr_RNIV7C99_S[16]\, 
        un3_rbinnext_cry_17, \rbinaddr_RNIJENN9_S[17]\, 
        un3_rbinnext_cry_18, \rbinaddr_RNI8M26A_S[18]\, 
        un3_rbinnext_cry_19, \rbinaddr_RNIUUDKA_S[19]\, 
        un3_rbinnext_cry_20, \rbinaddr_RNIC0Q2B_S[20]\, 
        un3_rbinnext_cry_21, \rbinaddr_RNIR26HB_S[21]\, 
        un3_rbinnext_cry_22, \rbinaddr_RNIB6IVB_S[22]\, 
        un3_rbinnext_cry_23, \rbinaddr_RNISAUDC_S[23]\, 
        un3_rbinnext_cry_24, \rbinaddr_RNIEGASC_S[24]\, 
        un3_rbinnext_cry_25, \rbinaddr_RNI1NMAD_S[25]\, 
        un3_rbinnext_cry_26, \rbinaddr_RNILU2PD_S[26]\, 
        un3_rbinnext_cry_27, \rbinaddr_RNIA7F7E_S[27]\, 
        un3_rbinnext_cry_28, \rbinaddr_RNI0HRLE_S[28]\, 
        un3_rbinnext_cry_29, \rbinaddr_RNINR74F_S[29]\, 
        un3_rbinnext_cry_30, \rbinaddr_RNI6VKIF_S[30]\, 
        un3_rbinnext_cry_31, \rbinaddr_RNIM321G_S[31]\, 
        un6_wbinnext_cry_0_cy, un6_wbinnext_cry_0, 
        \wbinaddr_RNIJ3OU_S[0]\, un6_wbinnext_cry_1, 
        \wbinaddr_RNIL3PD1_S[1]\, un6_wbinnext_cry_2, 
        \wbinaddr_RNIO4QS1_S[2]\, un6_wbinnext_cry_3, 
        \wbinaddr_RNIS6RB2_S[3]\, un6_wbinnext_cry_4, 
        \wbinaddr_RNI1ASQ2_S[4]\, un6_wbinnext_cry_5, 
        \wbinaddr_RNI7ET93_S[5]\, un6_wbinnext_cry_6, 
        \wbinaddr_RNIEJUO3_S[6]\, un6_wbinnext_cry_7, 
        \wbinaddr_RNIMPV74_S[7]\, un6_wbinnext_cry_8, 
        \wbinaddr_RNIV01N4_S[8]\, un6_wbinnext_cry_9, 
        \wbinaddr_RNI99265_S[9]\, un6_wbinnext_cry_10, 
        \wbinaddr_RNIRV1M5_S[10]\, un6_wbinnext_cry_11, 
        \wbinaddr_RNIEN166_S[11]\, un6_wbinnext_cry_12, 
        \wbinaddr_RNI2G1M6_S[12]\, un6_wbinnext_cry_13, 
        \wbinaddr_RNIN9167_S[13]\, un6_wbinnext_cry_14, 
        \wbinaddr_RNID41M7_S[14]\, un6_wbinnext_cry_15, 
        \wbinaddr_RNI40168_S[15]\, un6_wbinnext_cry_16, 
        \wbinaddr_RNISS0M8_S[16]\, un6_wbinnext_cry_17, 
        \wbinaddr_RNILQ069_S[17]\, un6_wbinnext_cry_18, 
        \wbinaddr_RNIFP0M9_S[18]\, un6_wbinnext_cry_19, 
        \wbinaddr_RNIAP06A_S[19]\, un6_wbinnext_cry_20, 
        \wbinaddr_RNITH16A_S[20]\, un6_wbinnext_cry_21, 
        \wbinaddr_RNIHB26A_S[21]\, un6_wbinnext_cry_22, 
        \wbinaddr_RNI6636A_S[22]\, un6_wbinnext_cry_23, 
        \wbinaddr_RNIS146A_S[23]\, un6_wbinnext_cry_24, 
        \wbinaddr_RNIJU46A_S[24]\, un6_wbinnext_cry_25, 
        \wbinaddr_RNIBS56A_S[25]\, un6_wbinnext_cry_26, 
        \wbinaddr_RNI4R66A_S[26]\, un6_wbinnext_cry_27, 
        \wbinaddr_RNIUQ76A_S[27]\, un6_wbinnext_cry_28, 
        \wbinaddr_RNIPR86A_S[28]\, un6_wbinnext_cry_29, 
        \wbinaddr_RNILT96A_S[29]\, un6_wbinnext_cry_30, 
        \wbinaddr_RNI9OB6A_S[30]\, un6_wbinnext_cry_31, 
        \wbinaddr_RNIUJD6A_S[31]\, 
        \fifo_empty_xhdl3_0_data_tmp[0]\, 
        fifo_empty_xhdl3_0_I_5_0, 
        \fifo_empty_xhdl3_0_data_tmp[1]\, 
        fifo_empty_xhdl3_0_I_77_0, 
        \fifo_empty_xhdl3_0_data_tmp[2]\, 
        fifo_empty_xhdl3_0_I_95_0, 
        \fifo_empty_xhdl3_0_data_tmp[3]\, 
        fifo_empty_xhdl3_0_I_89_0, 
        \fifo_empty_xhdl3_0_data_tmp[4]\, 
        fifo_empty_xhdl3_0_I_83_0, 
        \fifo_empty_xhdl3_0_data_tmp[5]\, 
        fifo_empty_xhdl3_0_I_53_0, 
        \fifo_empty_xhdl3_0_data_tmp[6]\, 
        fifo_empty_xhdl3_0_I_41_0, 
        \fifo_empty_xhdl3_0_data_tmp[7]\, 
        fifo_empty_xhdl3_0_I_47_0, 
        \fifo_empty_xhdl3_0_data_tmp[8]\, 
        fifo_empty_xhdl3_0_I_59_0, 
        \fifo_empty_xhdl3_0_data_tmp[9]\, 
        fifo_empty_xhdl3_0_I_29_0, 
        \fifo_empty_xhdl3_0_data_tmp[10]\, 
        fifo_empty_xhdl3_0_I_65_0, 
        \fifo_empty_xhdl3_0_data_tmp[11]\, 
        fifo_empty_xhdl3_0_I_71_0, 
        \fifo_empty_xhdl3_0_data_tmp[12]\, 
        fifo_empty_xhdl3_0_I_35_0, 
        \fifo_empty_xhdl3_0_data_tmp[13]\, 
        fifo_empty_xhdl3_0_I_23_0, 
        \fifo_empty_xhdl3_0_data_tmp[14]\, 
        fifo_empty_xhdl3_0_I_17_0, 
        \fifo_empty_xhdl3_0_data_tmp[15]\, 
        fifo_empty_xhdl3_0_I_11_0, \un13_writefull_0_data_tmp[0]\, 
        \un13_writefull_0_data_tmp[1]\, 
        \un13_writefull_0_data_tmp[2]\, 
        \un13_writefull_0_data_tmp[3]\, 
        \un13_writefull_0_data_tmp[4]\, 
        \un13_writefull_0_data_tmp[5]\, 
        \un13_writefull_0_data_tmp[6]\, 
        \un13_writefull_0_data_tmp[7]\, 
        \un13_writefull_0_data_tmp[8]\, 
        \un13_writefull_0_data_tmp[9]\, 
        \un13_writefull_0_data_tmp[10]\, un13_writefull_0_N_27, 
        \un13_writefull_0_data_tmp[11]\, 
        \un13_writefull_0_data_tmp[12]\, 
        \un13_writefull_0_data_tmp[13]\, 
        \un13_writefull_0_data_tmp[14]\, un13_writefull_0_N_2, 
        \un7_writefull\ : std_logic;

    for all : CoreAHBLtoAXI_wrch_ramHX
	Use entity work.CoreAHBLtoAXI_wrch_ramHX(DEF_ARCH);
begin 


    \wgraynext[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI99265_S[9]\, B => 
        \wbinaddr_RNIV01N4_S[8]\, Y => \wgraynext[8]_net_1\);
    
    \rbinaddr_RNI1H8L2[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_1, S
         => \rbinaddr_RNI1H8L2_S[2]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_2);
    
    \wgraynext[17]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIFP0M9_S[18]\, B => 
        \wbinaddr_RNILQ069_S[17]\, Y => \wgraynext[17]_net_1\);
    
    \wbinaddr_RNIEN166[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_10, S
         => \wbinaddr_RNIEN166_S[11]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_11);
    
    \Read_Bin_Ptr.rbinaddr_3[27]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIA7F7E_S[27]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[27]\);
    
    \raddr_gray[17]\ : SLE
      port map(D => \rgraynext[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[17]_net_1\);
    
    \rgraynext[28]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNINR74F_S[29]\, B => 
        \rbinaddr_RNI0HRLE_S[28]\, Y => \rgraynext[28]_net_1\);
    
    \rddata_r[55]\ : SLE
      port map(D => \port_xhdl7[55]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[55]_net_1\);
    
    \wgraynext[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIO4QS1_S[2]\, B => 
        \wbinaddr_RNIS6RB2_S[3]\, Y => \wgraynext[2]_net_1\);
    
    fifo_full_xhdl2_RNII4NF : ARI1
      generic map(INIT => x"40400")

      port map(A => wrch_fifo_wr_en_r, B => \fifo_full_xhdl2\, C
         => \wren_2\, D => ahb_busyidle_cyc, FCI => VCC_net_1, S
         => OPEN, Y => OPEN, FCO => un6_wbinnext_cry_0_cy);
    
    \Write_Bin_Ptr.wbinaddr_2[13]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIN9167_S[13]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[13]\);
    
    \rddata_r[23]\ : SLE
      port map(D => \port_xhdl7[23]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[23]_net_1\);
    
    \rddata_r_RNI3B0O[46]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[46]\, C => 
        \rddata_r[46]_net_1\, Y => N_288);
    
    \wsync2_rptr[2]\ : SLE
      port map(D => \wsync1_rptr[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[2]_net_1\);
    
    fifo_empty_xhdl3_RNO : CFG1
      generic map(INIT => "01")

      port map(A => fifo_empty_xhdl3_0_N_2, Y => 
        fifo_empty_xhdl3_0_N_2_i);
    
    \rsync2_wptr[30]\ : SLE
      port map(D => \rsync1_wptr[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[30]_net_1\);
    
    \rbinaddr[17]\ : SLE
      port map(D => \rbinaddr_3[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[17]_net_1\);
    
    \wbinaddr[4]\ : SLE
      port map(D => \wbinaddr_2[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[4]_net_1\);
    
    un13_writefull_0_I_51 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[17]_net_1\, B => 
        \wgraynext[16]_net_1\, C => \wgraynext[17]_net_1\, D => 
        \wsync2_rptr[16]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[7]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[8]\);
    
    \wsync2_rptr[0]\ : SLE
      port map(D => \wsync1_rptr[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[0]_net_1\);
    
    \rddata_r[34]\ : SLE
      port map(D => \port_xhdl7[34]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[34]_net_1\);
    
    \wgraynext[24]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIBS56A_S[25]\, B => 
        \wbinaddr_RNIJU46A_S[24]\, Y => \wgraynext[24]_net_1\);
    
    \rddata_r[61]\ : SLE
      port map(D => \port_xhdl7[61]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[61]_net_1\);
    
    \raddr_gray[14]\ : SLE
      port map(D => \rgraynext[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[14]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_39\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[13]_net_1\, B => 
        \rbinaddr_RNI9QAU7_S[13]\, C => \rbinaddr_RNIQTLC8_S[14]\, 
        D => fifo_empty_xhdl3_0_I_41_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[5]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[6]\);
    
    \rddata_r_RNI96851[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[2]\, C => 
        \rddata_r[2]_net_1\, Y => N_149);
    
    \rddata_r[58]\ : SLE
      port map(D => \port_xhdl7[58]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[58]_net_1\);
    
    \raddr_gray[31]\ : SLE
      port map(D => \rgraynext[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[31]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_29_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI8M26A_S[18]\, B => 
        \rsync2_wptr[18]_net_1\, Y => fifo_empty_xhdl3_0_I_29_0);
    
    \raddr_gray[16]\ : SLE
      port map(D => \rgraynext[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[16]_net_1\);
    
    \rddata_r[60]\ : SLE
      port map(D => \port_xhdl7[60]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[60]_net_1\);
    
    \rddata_r[25]\ : SLE
      port map(D => \port_xhdl7[25]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[25]_net_1\);
    
    un13_writefull_0_I_75 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[25]_net_1\, B => 
        \wgraynext[24]_net_1\, C => \wgraynext[25]_net_1\, D => 
        \wsync2_rptr[24]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[11]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[12]\);
    
    \rddata_r_RNI080O[43]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[43]\, C => 
        \rddata_r[43]_net_1\, Y => N_291);
    
    \Read_Bin_Ptr.rbinaddr_3[14]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIQTLC8_S[14]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[14]\);
    
    \rddata_r_RNIVNIU[16]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[16]\, C => 
        \rddata_r[16]_net_1\, Y => N_422);
    
    \rgraynext[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI32A52_S[1]\, B => 
        \rbinaddr_RNI6KBL1_S[0]\, Y => \rgraynext[0]_net_1\);
    
    un13_writefull_0_I_9 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[3]_net_1\, B => 
        \wgraynext[2]_net_1\, C => \wgraynext[3]_net_1\, D => 
        \wsync2_rptr[2]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[0]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[1]\);
    
    un13_writefull_0_I_27 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[9]_net_1\, B => 
        \wgraynext[8]_net_1\, C => \wgraynext[9]_net_1\, D => 
        \wsync2_rptr[8]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[3]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[4]\);
    
    \wgraynext[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI9OB6A_S[30]\, B => 
        \wbinaddr_RNILT96A_S[29]\, Y => \wgraynext[29]_net_1\);
    
    U_WRCH_RAM : CoreAHBLtoAXI_wrch_ramHX
      port map(port_xhdl7(63) => \port_xhdl7[63]\, port_xhdl7(62)
         => \port_xhdl7[62]\, port_xhdl7(61) => \port_xhdl7[61]\, 
        port_xhdl7(60) => \port_xhdl7[60]\, port_xhdl7(59) => 
        \port_xhdl7[59]\, port_xhdl7(58) => \port_xhdl7[58]\, 
        port_xhdl7(57) => \port_xhdl7[57]\, port_xhdl7(56) => 
        \port_xhdl7[56]\, port_xhdl7(55) => \port_xhdl7[55]\, 
        port_xhdl7(54) => \port_xhdl7[54]\, port_xhdl7(53) => 
        \port_xhdl7[53]\, port_xhdl7(52) => \port_xhdl7[52]\, 
        port_xhdl7(51) => \port_xhdl7[51]\, port_xhdl7(50) => 
        \port_xhdl7[50]\, port_xhdl7(49) => \port_xhdl7[49]\, 
        port_xhdl7(48) => \port_xhdl7[48]\, port_xhdl7(47) => 
        \port_xhdl7[47]\, port_xhdl7(46) => \port_xhdl7[46]\, 
        port_xhdl7(45) => \port_xhdl7[45]\, port_xhdl7(44) => 
        \port_xhdl7[44]\, port_xhdl7(43) => \port_xhdl7[43]\, 
        port_xhdl7(42) => \port_xhdl7[42]\, port_xhdl7(41) => 
        \port_xhdl7[41]\, port_xhdl7(40) => \port_xhdl7[40]\, 
        port_xhdl7(39) => \port_xhdl7[39]\, port_xhdl7(38) => 
        \port_xhdl7[38]\, port_xhdl7(37) => \port_xhdl7[37]\, 
        port_xhdl7(36) => \port_xhdl7[36]\, port_xhdl7(35) => 
        \port_xhdl7[35]\, port_xhdl7(34) => \port_xhdl7[34]\, 
        port_xhdl7(33) => \port_xhdl7[33]\, port_xhdl7(32) => 
        \port_xhdl7[32]\, port_xhdl7(31) => \port_xhdl7[31]\, 
        port_xhdl7(30) => \port_xhdl7[30]\, port_xhdl7(29) => 
        \port_xhdl7[29]\, port_xhdl7(28) => \port_xhdl7[28]\, 
        port_xhdl7(27) => \port_xhdl7[27]\, port_xhdl7(26) => 
        \port_xhdl7[26]\, port_xhdl7(25) => \port_xhdl7[25]\, 
        port_xhdl7(24) => \port_xhdl7[24]\, port_xhdl7(23) => 
        \port_xhdl7[23]\, port_xhdl7(22) => \port_xhdl7[22]\, 
        port_xhdl7(21) => \port_xhdl7[21]\, port_xhdl7(20) => 
        \port_xhdl7[20]\, port_xhdl7(19) => \port_xhdl7[19]\, 
        port_xhdl7(18) => \port_xhdl7[18]\, port_xhdl7(17) => 
        \port_xhdl7[17]\, port_xhdl7(16) => \port_xhdl7[16]\, 
        port_xhdl7(15) => \port_xhdl7[15]\, port_xhdl7(14) => 
        \port_xhdl7[14]\, port_xhdl7(13) => \port_xhdl7[13]\, 
        port_xhdl7(12) => \port_xhdl7[12]\, port_xhdl7(11) => 
        \port_xhdl7[11]\, port_xhdl7(10) => \port_xhdl7[10]\, 
        port_xhdl7(9) => \port_xhdl7[9]\, port_xhdl7(8) => 
        \port_xhdl7[8]\, port_xhdl7(7) => \port_xhdl7[7]\, 
        port_xhdl7(6) => \port_xhdl7[6]\, port_xhdl7(5) => 
        \port_xhdl7[5]\, port_xhdl7(4) => \port_xhdl7[4]\, 
        port_xhdl7(3) => \port_xhdl7[3]\, port_xhdl7(2) => 
        \port_xhdl7[2]\, port_xhdl7(1) => \port_xhdl7[1]\, 
        port_xhdl7(0) => \port_xhdl7[0]\, wrch_hwdata_r(31) => 
        wrch_hwdata_r(31), wrch_hwdata_r(30) => wrch_hwdata_r(30), 
        wrch_hwdata_r(29) => wrch_hwdata_r(29), wrch_hwdata_r(28)
         => wrch_hwdata_r(28), wrch_hwdata_r(27) => 
        wrch_hwdata_r(27), wrch_hwdata_r(26) => wrch_hwdata_r(26), 
        wrch_hwdata_r(25) => wrch_hwdata_r(25), wrch_hwdata_r(24)
         => wrch_hwdata_r(24), wrch_hwdata_r(23) => 
        wrch_hwdata_r(23), wrch_hwdata_r(22) => wrch_hwdata_r(22), 
        wrch_hwdata_r(21) => wrch_hwdata_r(21), wrch_hwdata_r(20)
         => wrch_hwdata_r(20), wrch_hwdata_r(19) => 
        wrch_hwdata_r(19), wrch_hwdata_r(18) => wrch_hwdata_r(18), 
        wrch_hwdata_r(17) => wrch_hwdata_r(17), wrch_hwdata_r(16)
         => wrch_hwdata_r(16), wrch_hwdata_r(15) => 
        wrch_hwdata_r(15), wrch_hwdata_r(14) => wrch_hwdata_r(14), 
        wrch_hwdata_r(13) => wrch_hwdata_r(13), wrch_hwdata_r(12)
         => wrch_hwdata_r(12), wrch_hwdata_r(11) => 
        wrch_hwdata_r(11), wrch_hwdata_r(10) => wrch_hwdata_r(10), 
        wrch_hwdata_r(9) => wrch_hwdata_r(9), wrch_hwdata_r(8)
         => wrch_hwdata_r(8), wrch_hwdata_r(7) => 
        wrch_hwdata_r(7), wrch_hwdata_r(6) => wrch_hwdata_r(6), 
        wrch_hwdata_r(5) => wrch_hwdata_r(5), wrch_hwdata_r(4)
         => wrch_hwdata_r(4), wrch_hwdata_r(3) => 
        wrch_hwdata_r(3), wrch_hwdata_r(2) => wrch_hwdata_r(2), 
        wrch_hwdata_r(1) => wrch_hwdata_r(1), wrch_hwdata_r(0)
         => wrch_hwdata_r(0), wbinaddr(3) => \wbinaddr[3]_net_1\, 
        wbinaddr(2) => \wbinaddr[2]_net_1\, wbinaddr(1) => 
        \wbinaddr[1]_net_1\, wbinaddr(0) => \wbinaddr[0]_net_1\, 
        rbinaddr(3) => \rbinaddr[3]_net_1\, rbinaddr(2) => 
        \rbinaddr[2]_net_1\, rbinaddr(1) => \rbinaddr[1]_net_1\, 
        rbinaddr(0) => \rbinaddr[0]_net_1\, wrch_fifo_wr_en_r => 
        wrch_fifo_wr_en_r, fifo_full_xhdl2 => \fifo_full_xhdl2\, 
        wren_2 => \wren_2\, SDRCLK_c => SDRCLK_c);
    
    \Read_Bin_Ptr.rbinaddr_3[26]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNILU2PD_S[26]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[26]\);
    
    \Read_Bin_Ptr.rbinaddr_3[11]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIAMK17_S[11]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[11]\);
    
    \rddata_r_RNIB8851[4]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[4]\, C => 
        \rddata_r[4]_net_1\, Y => N_147);
    
    \rddata_r[28]\ : SLE
      port map(D => \port_xhdl7[28]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[28]_net_1\);
    
    \rbinaddr_RNI01753[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_2, S
         => \rbinaddr_RNI01753_S[3]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_3);
    
    \rddata_r[54]\ : SLE
      port map(D => \port_xhdl7[54]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[54]_net_1\);
    
    un13_writefull_0_I_39 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[13]_net_1\, B => 
        \wgraynext[12]_net_1\, C => \wgraynext[13]_net_1\, D => 
        \wsync2_rptr[12]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[5]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[6]\);
    
    \wbinaddr[18]\ : SLE
      port map(D => \wbinaddr_2[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[18]_net_1\);
    
    \rddata_r_RNI0QJU[26]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[26]\, C => 
        \rddata_r[26]_net_1\, Y => N_417);
    
    \rgraynext[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIPNVF7_S[12]\, B => 
        \rbinaddr_RNIAMK17_S[11]\, Y => \rgraynext[11]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[18]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIFP0M9_S[18]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[18]\);
    
    \wbinaddr[19]\ : SLE
      port map(D => \wbinaddr_2[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[19]_net_1\);
    
    \rbinaddr[25]\ : SLE
      port map(D => \rbinaddr_3[25]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[25]_net_1\);
    
    \raddr_gray[2]\ : SLE
      port map(D => \rgraynext[2]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[2]_net_1\);
    
    \wbinaddr[27]\ : SLE
      port map(D => \wbinaddr_2[27]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[27]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[22]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI6636A_S[22]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[22]\);
    
    \rsync2_wptr[8]\ : SLE
      port map(D => \rsync1_wptr[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[8]_net_1\);
    
    \rgraynext[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0I5L3_S[4]\, B => 
        \rbinaddr_RNI01753_S[3]\, Y => \rgraynext[3]_net_1\);
    
    \wbinaddr_RNILT96A[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_28, S
         => \wbinaddr_RNILT96A_S[29]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_29);
    
    \rsync1_wptr[12]\ : SLE
      port map(D => \waddr_gray[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[12]_net_1\);
    
    \rgraynext[26]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIA7F7E_S[27]\, B => 
        \rbinaddr_RNILU2PD_S[26]\, Y => \rgraynext[26]_net_1\);
    
    \rsync2_wptr[12]\ : SLE
      port map(D => \rsync1_wptr[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[12]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_89_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI3N2L4_S[6]\, B => 
        \rsync2_wptr[6]_net_1\, Y => fifo_empty_xhdl3_0_I_89_0);
    
    \rddata_r_RNIDA851[6]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[6]\, C => 
        \rddata_r[6]_net_1\, Y => N_411);
    
    \rbinaddr[21]\ : SLE
      port map(D => \rbinaddr_3[21]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[21]_net_1\);
    
    \wsync2_rptr[8]\ : SLE
      port map(D => \wsync1_rptr[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[8]_net_1\);
    
    \rddata_r[24]\ : SLE
      port map(D => \port_xhdl7[24]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[24]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_47_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIQTLC8_S[14]\, B => 
        \rsync2_wptr[14]_net_1\, Y => fifo_empty_xhdl3_0_I_47_0);
    
    \rgraynext[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIFMU46_S[9]\, B => 
        \rbinaddr_RNIA00L5_S[8]\, Y => \rgraynext[8]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[20]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIC0Q2B_S[20]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[20]\);
    
    \rddata_r_RNIV5VN[33]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[33]\, C => 
        \rddata_r[33]_net_1\, Y => N_159);
    
    \wgraynext[23]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIJU46A_S[24]\, B => 
        \wbinaddr_RNIS146A_S[23]\, Y => \wgraynext[23]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_27\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[19]_net_1\, B => 
        \rbinaddr_RNIUUDKA_S[19]\, C => \rbinaddr_RNIC0Q2B_S[20]\, 
        D => fifo_empty_xhdl3_0_I_29_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[8]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[9]\);
    
    \waddr_gray[11]\ : SLE
      port map(D => \wgraynext[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[11]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[1]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI32A52_S[1]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[1]\);
    
    \Read_Bin_Ptr.rbinaddr_3[15]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIC21R8_S[15]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[15]\);
    
    \wgraynext[22]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIS146A_S[23]\, B => 
        \wbinaddr_RNI6636A_S[22]\, Y => \wgraynext[22]_net_1\);
    
    \waddr_gray[26]\ : SLE
      port map(D => \wgraynext[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[26]_net_1\);
    
    \rddata_r[42]\ : SLE
      port map(D => \port_xhdl7[42]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[42]_net_1\);
    
    \rgraynext[17]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI8M26A_S[18]\, B => 
        \rbinaddr_RNIJENN9_S[17]\, Y => \rgraynext[17]_net_1\);
    
    \rddata_r_RNI2A0O[45]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[45]\, C => 
        \rddata_r[45]_net_1\, Y => N_289);
    
    \Write_Bin_Ptr.wbinaddr_2[31]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIUJD6A_S[31]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[31]\);
    
    \rsync1_wptr[2]\ : SLE
      port map(D => \waddr_gray[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[2]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_5_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI6KBL1_S[0]\, B => 
        \rsync2_wptr[0]_net_1\, Y => fifo_empty_xhdl3_0_I_5_0);
    
    \rgraynext[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI14454_S[5]\, B => 
        \rbinaddr_RNI0I5L3_S[4]\, Y => \rgraynext[4]_net_1\);
    
    \rgraynext[25]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNILU2PD_S[26]\, B => 
        \rbinaddr_RNI1NMAD_S[25]\, Y => \rgraynext[25]_net_1\);
    
    \rddata_r[13]\ : SLE
      port map(D => \port_xhdl7[13]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[13]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_33\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[25]_net_1\, B => 
        \rbinaddr_RNI1NMAD_S[25]\, C => \rbinaddr_RNILU2PD_S[26]\, 
        D => fifo_empty_xhdl3_0_I_35_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[11]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[12]\);
    
    \waddr_gray[10]\ : SLE
      port map(D => \wgraynext[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[10]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_15\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[29]_net_1\, B => 
        \rbinaddr_RNINR74F_S[29]\, C => \rbinaddr_RNI6VKIF_S[30]\, 
        D => fifo_empty_xhdl3_0_I_17_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[13]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[14]\);
    
    \rddata_r_RNIQJJU[20]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[20]\, C => 
        \rddata_r[20]_net_1\, Y => N_214);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_23_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNILU2PD_S[26]\, B => 
        \rsync2_wptr[26]_net_1\, Y => fifo_empty_xhdl3_0_I_23_0);
    
    \rddata_r_RNI2B2O[62]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[62]\, C => 
        \rddata_r[62]_net_1\, Y => N_328);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_9\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[31]_net_1\, B => 
        \rbinaddr_RNIM321G_S[31]\, C => \rbinaddr_RNI79FFG_S[32]\, 
        D => fifo_empty_xhdl3_0_I_11_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[14]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[15]\);
    
    \rsync2_wptr[6]\ : SLE
      port map(D => \rsync1_wptr[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[6]_net_1\);
    
    \rsync1_wptr[25]\ : SLE
      port map(D => \waddr_gray[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[25]_net_1\);
    
    \waddr_gray[8]\ : SLE
      port map(D => \wgraynext[8]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[8]_net_1\);
    
    \rbinaddr_RNIB6IVB[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_21, S
         => \rbinaddr_RNIB6IVB_S[22]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_22);
    
    \wsync2_rptr[28]\ : SLE
      port map(D => \wsync1_rptr[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[28]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_35_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIEGASC_S[24]\, B => 
        \rsync2_wptr[24]_net_1\, Y => fifo_empty_xhdl3_0_I_35_0);
    
    \rbinaddr[24]\ : SLE
      port map(D => \rbinaddr_3[24]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[24]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[6]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIEJUO3_S[6]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[6]\);
    
    \wgraynext[18]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIAP06A_S[19]\, B => 
        \wbinaddr_RNIFP0M9_S[18]\, Y => \wgraynext[18]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[2]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI1H8L2_S[2]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[2]\);
    
    \wbinaddr[22]\ : SLE
      port map(D => \wbinaddr_2[22]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[22]_net_1\);
    
    \wsync2_rptr[18]\ : SLE
      port map(D => \wsync1_rptr[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[18]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_69\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[23]_net_1\, B => 
        \rbinaddr_RNISAUDC_S[23]\, C => \rbinaddr_RNIEGASC_S[24]\, 
        D => fifo_empty_xhdl3_0_I_71_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[10]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[11]\);
    
    \rddata_r[15]\ : SLE
      port map(D => \port_xhdl7[15]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[15]_net_1\);
    
    \wgraynext[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIV01N4_S[8]\, B => 
        \wbinaddr_RNIMPV74_S[7]\, Y => \wgraynext[7]_net_1\);
    
    \wgraynext[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI7ET93_S[5]\, B => 
        \wbinaddr_RNI1ASQ2_S[4]\, Y => \wgraynext[4]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \rgraynext[24]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI1NMAD_S[25]\, B => 
        \rbinaddr_RNIEGASC_S[24]\, Y => \rgraynext[24]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[14]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNID41M7_S[14]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[14]\);
    
    \rddata_r_RNI5D1O[56]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[56]\, C => 
        \rddata_r[56]_net_1\, Y => N_421);
    
    \rbinaddr[23]\ : SLE
      port map(D => \rbinaddr_3[23]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[23]_net_1\);
    
    \rsync2_wptr[29]\ : SLE
      port map(D => \rsync1_wptr[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[29]_net_1\);
    
    un13_writefull_0_I_45 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[15]_net_1\, B => 
        \wgraynext[14]_net_1\, C => \wgraynext[15]_net_1\, D => 
        \wsync2_rptr[14]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[6]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[7]\);
    
    \rbinaddr[26]\ : SLE
      port map(D => \rbinaddr_3[26]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[26]_net_1\);
    
    \rddata_r_RNISLJU[22]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[22]\, C => 
        \rddata_r[22]_net_1\, Y => N_436);
    
    \raddr_gray[10]\ : SLE
      port map(D => \rgraynext[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[10]_net_1\);
    
    \raddr_gray[25]\ : SLE
      port map(D => \rgraynext[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[25]_net_1\);
    
    \waddr_gray[13]\ : SLE
      port map(D => \wgraynext[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[13]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[23]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNISAUDC_S[23]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[23]\);
    
    \wbinaddr[20]\ : SLE
      port map(D => \wbinaddr_2[20]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[20]_net_1\);
    
    \rbinaddr[1]\ : SLE
      port map(D => \rbinaddr_3[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[1]_net_1\);
    
    \rddata_r[18]\ : SLE
      port map(D => \port_xhdl7[18]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[18]_net_1\);
    
    \raddr_gray[28]\ : SLE
      port map(D => \rgraynext[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[28]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[11]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIEN166_S[11]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[11]\);
    
    \wsync2_rptr[32]\ : SLE
      port map(D => \wsync1_rptr[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[32]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[2]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIO4QS1_S[2]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[2]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_83_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIA00L5_S[8]\, B => 
        \rsync2_wptr[8]_net_1\, Y => fifo_empty_xhdl3_0_I_83_0);
    
    \rddata_r[32]\ : SLE
      port map(D => \port_xhdl7[32]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[32]_net_1\);
    
    \rgraynext[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI6VKIF_S[30]\, B => 
        \rbinaddr_RNINR74F_S[29]\, Y => \rgraynext[29]_net_1\);
    
    \wbinaddr[25]\ : SLE
      port map(D => \wbinaddr_2[25]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[25]_net_1\);
    
    \rbinaddr[15]\ : SLE
      port map(D => \rbinaddr_3[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[15]_net_1\);
    
    \wbinaddr[17]\ : SLE
      port map(D => \wbinaddr_2[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[17]_net_1\);
    
    \waddr_gray[9]\ : SLE
      port map(D => \wgraynext[9]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[9]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[0]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIJ3OU_S[0]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[0]\);
    
    \rddata_r_RNIRKIU[13]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[13]\, C => 
        \rddata_r[13]_net_1\, Y => N_282);
    
    \rddata_r_RNIV60O[42]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[42]\, C => 
        \rddata_r[42]_net_1\, Y => N_292);
    
    \rddata_r_RNI18VN[35]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[35]\, C => 
        \rddata_r[35]_net_1\, Y => N_157);
    
    \rbinaddr[11]\ : SLE
      port map(D => \rbinaddr_3[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[11]_net_1\);
    
    \rsync1_wptr[4]\ : SLE
      port map(D => \waddr_gray[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[4]_net_1\);
    
    \rsync1_wptr[32]\ : SLE
      port map(D => \waddr_gray[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[32]_net_1\);
    
    \rddata_r[63]\ : SLE
      port map(D => \port_xhdl7[63]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[63]_net_1\);
    
    \rsync2_wptr[32]\ : SLE
      port map(D => \rsync1_wptr[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[32]_net_1\);
    
    \waddr_gray[29]\ : SLE
      port map(D => \wgraynext[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[29]_net_1\);
    
    \rddata_r[14]\ : SLE
      port map(D => \port_xhdl7[14]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[14]_net_1\);
    
    \rbinaddr[8]\ : SLE
      port map(D => \rbinaddr_3[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[8]_net_1\);
    
    \wbinaddr_RNI4R66A[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_25, S
         => \wbinaddr_RNI4R66A_S[26]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_26);
    
    \rddata_r[52]\ : SLE
      port map(D => \port_xhdl7[52]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[52]_net_1\);
    
    \wbinaddr_RNIMPV74[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_6, S
         => \wbinaddr_RNIMPV74_S[7]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_7);
    
    \rbinaddr_RNIC0Q2B[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_19, S
         => \rbinaddr_RNIC0Q2B_S[20]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_20);
    
    \rddata_r[7]\ : SLE
      port map(D => \port_xhdl7[7]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[7]_net_1\);
    
    \raddr_gray[27]\ : SLE
      port map(D => \rgraynext[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[27]_net_1\);
    
    \wsync1_rptr[22]\ : SLE
      port map(D => \raddr_gray[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[22]_net_1\);
    
    \wgraynext[16]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNILQ069_S[17]\, B => 
        \wbinaddr_RNISS0M8_S[16]\, Y => \wgraynext[16]_net_1\);
    
    \rgraynext[23]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIEGASC_S[24]\, B => 
        \rbinaddr_RNISAUDC_S[23]\, Y => \rgraynext[23]_net_1\);
    
    \rddata_r_RNI081O[51]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[51]\, C => 
        \rddata_r[51]_net_1\, Y => N_223);
    
    \rddata_r_RNI191O[52]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[52]\, C => 
        \rddata_r[52]_net_1\, Y => N_222);
    
    \rbinaddr_RNI6B155[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_6, S
         => \rbinaddr_RNI6B155_S[7]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_7);
    
    \Read_Bin_Ptr.rbinaddr_3[24]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIEGASC_S[24]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[24]\);
    
    \wsync1_rptr[21]\ : SLE
      port map(D => \raddr_gray[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[21]_net_1\);
    
    \rgraynext[22]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNISAUDC_S[23]\, B => 
        \rbinaddr_RNIB6IVB_S[22]\, Y => \rgraynext[22]_net_1\);
    
    \wsync1_rptr[12]\ : SLE
      port map(D => \raddr_gray[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[12]_net_1\);
    
    \rbinaddr_RNIFMU46[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_8, S
         => \rbinaddr_RNIFMU46_S[9]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_9);
    
    \rsync1_wptr[15]\ : SLE
      port map(D => \waddr_gray[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[15]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_21\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[27]_net_1\, B => 
        \rbinaddr_RNIA7F7E_S[27]\, C => \rbinaddr_RNI0HRLE_S[28]\, 
        D => fifo_empty_xhdl3_0_I_23_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[12]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[13]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_63\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[21]_net_1\, B => 
        \rbinaddr_RNIR26HB_S[21]\, C => \rbinaddr_RNIB6IVB_S[22]\, 
        D => fifo_empty_xhdl3_0_I_65_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[9]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[10]\);
    
    \wsync1_rptr[11]\ : SLE
      port map(D => \raddr_gray[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[11]_net_1\);
    
    \rddata_r_RNI1RJU[27]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[27]\, C => 
        \rddata_r[27]_net_1\, Y => N_438);
    
    \Read_Bin_Ptr.rbinaddr_3[21]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIR26HB_S[21]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[21]\);
    
    \raddr_gray[24]\ : SLE
      port map(D => \rgraynext[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[24]_net_1\);
    
    \rsync1_wptr[5]\ : SLE
      port map(D => \waddr_gray[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[5]_net_1\);
    
    \rddata_r[22]\ : SLE
      port map(D => \port_xhdl7[22]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[22]_net_1\);
    
    \rbinaddr[14]\ : SLE
      port map(D => \rbinaddr_3[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[14]_net_1\);
    
    \rgraynext[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIM321G_S[31]\, B => 
        \rbinaddr_RNI6VKIF_S[30]\, Y => \rgraynext[30]_net_1\);
    
    \rddata_r[49]\ : SLE
      port map(D => \port_xhdl7[49]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[49]_net_1\);
    
    \raddr_gray[26]\ : SLE
      port map(D => \rgraynext[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[26]_net_1\);
    
    \rgraynext[18]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIUUDKA_S[19]\, B => 
        \rbinaddr_RNI8M26A_S[18]\, Y => \rgraynext[18]_net_1\);
    
    \wbinaddr[12]\ : SLE
      port map(D => \wbinaddr_2[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[12]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[19]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIAP06A_S[19]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[19]\);
    
    \rbinaddr[31]\ : SLE
      port map(D => \rbinaddr_3[31]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[31]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[25]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIBS56A_S[25]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[25]\);
    
    \wbinaddr[21]\ : SLE
      port map(D => \wbinaddr_2[21]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[21]_net_1\);
    
    \rsync2_wptr[3]\ : SLE
      port map(D => \rsync1_wptr[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[3]_net_1\);
    
    \wgraynext[15]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNISS0M8_S[16]\, B => 
        \wbinaddr_RNI40168_S[15]\, Y => \wgraynext[15]_net_1\);
    
    \rsync2_wptr[19]\ : SLE
      port map(D => \rsync1_wptr[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[19]_net_1\);
    
    \rddata_r_RNI74851[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[0]\, C => 
        \rddata_r[0]_net_1\, Y => N_151);
    
    \rbinaddr[13]\ : SLE
      port map(D => \rbinaddr_3[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[13]_net_1\);
    
    \rddata_r_RNI1A2O[61]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[61]\, C => 
        \rddata_r[61]_net_1\, Y => N_432);
    
    \rddata_r[46]\ : SLE
      port map(D => \port_xhdl7[46]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[46]_net_1\);
    
    \rbinaddr[16]\ : SLE
      port map(D => \rbinaddr_3[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[16]_net_1\);
    
    un7_writefull : CFG2
      generic map(INIT => x"6")

      port map(A => \wgraynext[31]_net_1\, B => 
        \wsync2_rptr[31]_net_1\, Y => \un7_writefull\);
    
    \rddata_r_RNIC9851[5]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[5]\, C => 
        \rddata_r[5]_net_1\, Y => N_433);
    
    \wbinaddr[1]\ : SLE
      port map(D => \wbinaddr_2[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[1]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[20]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNITH16A_S[20]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[20]\);
    
    \rsync1_wptr[27]\ : SLE
      port map(D => \waddr_gray[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[27]_net_1\);
    
    \rbinaddr_RNINR74F[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_28, S
         => \rbinaddr_RNINR74F_S[29]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_29);
    
    \Write_Bin_Ptr.wbinaddr_2[4]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI1ASQ2_S[4]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[4]\);
    
    \wbinaddr[10]\ : SLE
      port map(D => \wbinaddr_2[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[10]_net_1\);
    
    \wbinaddr_RNIKGF6A[32]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[32]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_31, S
         => \wbinaddr_RNIKGF6A_S[32]\, Y => OPEN, FCO => OPEN);
    
    \wbinaddr_RNIV01N4[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_7, S
         => \wbinaddr_RNIV01N4_S[8]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_8);
    
    \wbinaddr_RNI99265[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_8, S
         => \wbinaddr_RNI99265_S[9]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_9);
    
    \wgraynext[14]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI40168_S[15]\, B => 
        \wbinaddr_RNID41M7_S[14]\, Y => \wgraynext[14]_net_1\);
    
    \wbinaddr[15]\ : SLE
      port map(D => \wbinaddr_2[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[15]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[25]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI1NMAD_S[25]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[25]\);
    
    \wbinaddr_RNIEJUO3[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_5, S
         => \wbinaddr_RNIEJUO3_S[6]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_6);
    
    \Read_Bin_Ptr.rbinaddr_3[9]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIFMU46_S[9]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[9]\);
    
    \waddr_gray[7]\ : SLE
      port map(D => \wgraynext[7]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[7]_net_1\);
    
    \rbinaddr[5]\ : SLE
      port map(D => \rbinaddr_3[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[5]_net_1\);
    
    \waddr_gray[14]\ : SLE
      port map(D => \wgraynext[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[14]_net_1\);
    
    \wbinaddr[32]\ : SLE
      port map(D => \wbinaddr_2[32]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[32]_net_1\);
    
    \raddr_gray[8]\ : SLE
      port map(D => \rgraynext[8]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[8]_net_1\);
    
    \wbinaddr[8]\ : SLE
      port map(D => \wbinaddr_2[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[8]_net_1\);
    
    \rddata_r_RNI29VN[36]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[36]\, C => 
        \rddata_r[36]_net_1\, Y => N_156);
    
    wren_1 : CFG2
      generic map(INIT => x"2")

      port map(A => wrch_fifo_wr_en_r, B => \wren_2\, Y => 
        \wren_1\);
    
    \rbinaddr_RNI8M26A[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_17, S
         => \rbinaddr_RNI8M26A_S[18]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_18);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_45\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[15]_net_1\, B => 
        \rbinaddr_RNIC21R8_S[15]\, C => \rbinaddr_RNIV7C99_S[16]\, 
        D => fifo_empty_xhdl3_0_I_47_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[6]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[7]\);
    
    \wsync1_rptr[1]\ : SLE
      port map(D => \raddr_gray[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[1]_net_1\);
    
    \waddr_gray[21]\ : SLE
      port map(D => \wgraynext[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[21]_net_1\);
    
    \wgraynext[19]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNITH16A_S[20]\, B => 
        \wbinaddr_RNIAP06A_S[19]\, Y => \wgraynext[19]_net_1\);
    
    \wbinaddr_RNIS146A[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_22, S
         => \wbinaddr_RNIS146A_S[23]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_23);
    
    \rddata_r[39]\ : SLE
      port map(D => \port_xhdl7[39]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[39]_net_1\);
    
    \waddr_gray[4]\ : SLE
      port map(D => \wgraynext[4]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[4]_net_1\);
    
    \rddata_r_RNI7E0O[49]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[49]\, C => 
        \rddata_r[49]_net_1\, Y => N_419);
    
    \rbinaddr[0]\ : SLE
      port map(D => \rbinaddr_3[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[0]_net_1\);
    
    \rsync2_wptr[28]\ : SLE
      port map(D => \rsync1_wptr[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[28]_net_1\);
    
    \rsync1_wptr[28]\ : SLE
      port map(D => \waddr_gray[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[28]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[3]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI01753_S[3]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[3]\);
    
    \rddata_r_RNIRLKU[30]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[30]\, C => 
        \rddata_r[30]_net_1\, Y => N_440);
    
    \wgraynext[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIMPV74_S[7]\, B => 
        \wbinaddr_RNIEJUO3_S[6]\, Y => \wgraynext[6]_net_1\);
    
    \rgraynext[16]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIJENN9_S[17]\, B => 
        \rbinaddr_RNIV7C99_S[16]\, Y => \rgraynext[16]_net_1\);
    
    \wgraynext[20]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIHB26A_S[21]\, B => 
        \wbinaddr_RNITH16A_S[20]\, Y => \wgraynext[20]_net_1\);
    
    \wbinaddr_RNIPR86A[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_27, S
         => \wbinaddr_RNIPR86A_S[28]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_28);
    
    \rddata_r[2]\ : SLE
      port map(D => \port_xhdl7[2]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[2]_net_1\);
    
    \wbinaddr[30]\ : SLE
      port map(D => \wbinaddr_2[30]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[30]_net_1\);
    
    \rddata_r[36]\ : SLE
      port map(D => \port_xhdl7[36]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[36]_net_1\);
    
    \waddr_gray[20]\ : SLE
      port map(D => \wgraynext[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[20]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[18]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI8M26A_S[18]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[18]\);
    
    \wgraynext[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIUJD6A_S[31]\, B => 
        \wbinaddr_RNI9OB6A_S[30]\, Y => \wgraynext[30]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[32]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIKGF6A_S[32]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[32]\);
    
    \wsync1_rptr[9]\ : SLE
      port map(D => \raddr_gray[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[9]_net_1\);
    
    \rddata_r[59]\ : SLE
      port map(D => \port_xhdl7[59]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[59]_net_1\);
    
    \rddata_r[12]\ : SLE
      port map(D => \port_xhdl7[12]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[12]_net_1\);
    
    \rsync1_wptr[7]\ : SLE
      port map(D => \waddr_gray[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[7]_net_1\);
    
    \raddr_gray[9]\ : SLE
      port map(D => \rgraynext[9]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[9]_net_1\);
    
    \wgraynext[13]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNID41M7_S[14]\, B => 
        \wbinaddr_RNIN9167_S[13]\, Y => \wgraynext[13]_net_1\);
    
    \wbinaddr[26]\ : SLE
      port map(D => \wbinaddr_2[26]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[26]_net_1\);
    
    \wbinaddr[11]\ : SLE
      port map(D => \wbinaddr_2[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[11]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[8]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIV01N4_S[8]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[8]\);
    
    \rgraynext[15]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIV7C99_S[16]\, B => 
        \rbinaddr_RNIC21R8_S[15]\, Y => \rgraynext[15]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_11_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI6VKIF_S[30]\, B => 
        \rsync2_wptr[30]_net_1\, Y => fifo_empty_xhdl3_0_I_11_0);
    
    \rddata_r_RNIU4VN[32]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[32]\, C => 
        \rddata_r[32]_net_1\, Y => N_160);
    
    un13_writefull_0_I_15 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[5]_net_1\, B => 
        \wgraynext[4]_net_1\, C => \wgraynext[5]_net_1\, D => 
        \wsync2_rptr[4]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[1]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[2]\);
    
    \wgraynext[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIN9167_S[13]\, B => 
        \wbinaddr_RNI2G1M6_S[12]\, Y => \wgraynext[12]_net_1\);
    
    \rddata_r[56]\ : SLE
      port map(D => \port_xhdl7[56]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[56]_net_1\);
    
    \rddata_r_RNI6D0O[48]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[48]\, C => 
        \rddata_r[48]_net_1\, Y => N_418);
    
    \wbinaddr_RNIS6RB2[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_2, S
         => \wbinaddr_RNIS6RB2_S[3]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_3);
    
    \raddr_gray[20]\ : SLE
      port map(D => \rgraynext[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[20]_net_1\);
    
    \raddr_gray[12]\ : SLE
      port map(D => \rgraynext[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[12]_net_1\);
    
    \wsync1_rptr[20]\ : SLE
      port map(D => \raddr_gray[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[20]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[7]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIMPV74_S[7]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[7]\);
    
    \rsync1_wptr[17]\ : SLE
      port map(D => \waddr_gray[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[17]_net_1\);
    
    \waddr_gray[23]\ : SLE
      port map(D => \wgraynext[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[23]_net_1\);
    
    \wsync1_rptr[26]\ : SLE
      port map(D => \raddr_gray[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[26]_net_1\);
    
    \rddata_r[29]\ : SLE
      port map(D => \port_xhdl7[29]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[29]_net_1\);
    
    \rsync1_wptr[21]\ : SLE
      port map(D => \waddr_gray[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[21]_net_1\);
    
    \rbinaddr[9]\ : SLE
      port map(D => \rbinaddr_3[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[9]_net_1\);
    
    \wsync1_rptr[10]\ : SLE
      port map(D => \raddr_gray[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[10]_net_1\);
    
    \rgraynext[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIA00L5_S[8]\, B => 
        \rbinaddr_RNI6B155_S[7]\, Y => \rgraynext[7]_net_1\);
    
    \rgraynext[14]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIC21R8_S[15]\, B => 
        \rbinaddr_RNIQTLC8_S[14]\, Y => \rgraynext[14]_net_1\);
    
    \wsync1_rptr[16]\ : SLE
      port map(D => \raddr_gray[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[16]_net_1\);
    
    \rddata_r[26]\ : SLE
      port map(D => \port_xhdl7[26]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[26]_net_1\);
    
    \wbinaddr[5]\ : SLE
      port map(D => \wbinaddr_2[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[5]_net_1\);
    
    \wsync2_rptr[20]\ : SLE
      port map(D => \wsync1_rptr[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[20]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[9]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI99265_S[9]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[9]\);
    
    \Write_Bin_Ptr.wbinaddr_2[12]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI2G1M6_S[12]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[12]\);
    
    \rddata_r_RNIRKJU[21]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[21]\, C => 
        \rddata_r[21]_net_1\, Y => N_213);
    
    \Write_Bin_Ptr.wbinaddr_2[26]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI4R66A_S[26]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[26]\);
    
    un13_writefull_0_I_57 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[19]_net_1\, B => 
        \wgraynext[18]_net_1\, C => \wgraynext[19]_net_1\, D => 
        \wsync2_rptr[18]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[8]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[9]\);
    
    \rsync1_wptr[24]\ : SLE
      port map(D => \waddr_gray[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[24]_net_1\);
    
    \wbinaddr[31]\ : SLE
      port map(D => \wbinaddr_2[31]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[31]_net_1\);
    
    \rbinaddr_RNIAMK17[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_10, S
         => \rbinaddr_RNIAMK17_S[11]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_11);
    
    \wsync2_rptr[10]\ : SLE
      port map(D => \wsync1_rptr[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[10]_net_1\);
    
    \wbinaddr[0]\ : SLE
      port map(D => \wbinaddr_2[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[0]_net_1\);
    
    \wgraynext[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIEJUO3_S[6]\, B => 
        \wbinaddr_RNI7ET93_S[5]\, Y => \wgraynext[5]_net_1\);
    
    \rgraynext[19]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIC0Q2B_S[20]\, B => 
        \rbinaddr_RNIUUDKA_S[19]\, Y => \rgraynext[19]_net_1\);
    
    \rddata_r_RNI5CVN[39]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[39]\, C => 
        \rddata_r[39]_net_1\, Y => N_427);
    
    \rsync2_wptr[26]\ : SLE
      port map(D => \rsync1_wptr[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[26]_net_1\);
    
    \wsync1_rptr[24]\ : SLE
      port map(D => \raddr_gray[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[24]_net_1\);
    
    \waddr_gray[17]\ : SLE
      port map(D => \wgraynext[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[17]_net_1\);
    
    \rsync2_wptr[18]\ : SLE
      port map(D => \rsync1_wptr[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[18]_net_1\);
    
    \rsync1_wptr[18]\ : SLE
      port map(D => \waddr_gray[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[18]_net_1\);
    
    \rddata_r_RNI8G1O[59]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[59]\, C => 
        \rddata_r[59]_net_1\, Y => N_431);
    
    \wsync2_rptr[1]\ : SLE
      port map(D => \wsync1_rptr[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[1]_net_1\);
    
    \wsync1_rptr[28]\ : SLE
      port map(D => \raddr_gray[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[28]_net_1\);
    
    \rddata_r[5]\ : SLE
      port map(D => \port_xhdl7[5]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[5]_net_1\);
    
    \rsync1_wptr[0]\ : SLE
      port map(D => \waddr_gray[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[0]_net_1\);
    
    \rddata_r[62]\ : SLE
      port map(D => \port_xhdl7[62]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[62]_net_1\);
    
    \wsync1_rptr[14]\ : SLE
      port map(D => \raddr_gray[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[14]_net_1\);
    
    \waddr_gray[31]\ : SLE
      port map(D => \wgraynext[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[31]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[3]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIS6RB2_S[3]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[3]\);
    
    \rbinaddr_RNIJENN9[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_16, S
         => \rbinaddr_RNIJENN9_S[17]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_17);
    
    \wsync1_rptr[18]\ : SLE
      port map(D => \raddr_gray[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[18]_net_1\);
    
    \wbinaddr_RNIRV1M5[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_9, S
         => \wbinaddr_RNIRV1M5_S[10]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_10);
    
    \rsync2_wptr[2]\ : SLE
      port map(D => \rsync1_wptr[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[2]_net_1\);
    
    \wbinaddr_RNI40168[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_14, S
         => \wbinaddr_RNI40168_S[15]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_15);
    
    \wsync1_rptr[23]\ : SLE
      port map(D => \raddr_gray[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[23]_net_1\);
    
    \rddata_r_RNI0PIU[17]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[17]\, C => 
        \rddata_r[17]_net_1\, Y => N_423);
    
    \rbinaddr[28]\ : SLE
      port map(D => \rbinaddr_3[28]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[28]_net_1\);
    
    \rddata_r[47]\ : SLE
      port map(D => \port_xhdl7[47]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[47]_net_1\);
    
    \wsync2_rptr[24]\ : SLE
      port map(D => \wsync1_rptr[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[24]_net_1\);
    
    \rgraynext[20]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIR26HB_S[21]\, B => 
        \rbinaddr_RNIC0Q2B_S[20]\, Y => \rgraynext[20]_net_1\);
    
    \waddr_gray[30]\ : SLE
      port map(D => \wgraynext[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[30]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[19]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIUUDKA_S[19]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[19]\);
    
    \wsync1_rptr[13]\ : SLE
      port map(D => \raddr_gray[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[13]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[27]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIUQ76A_S[27]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[27]\);
    
    \wsync2_rptr[9]\ : SLE
      port map(D => \wsync1_rptr[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[9]_net_1\);
    
    \wsync2_rptr[14]\ : SLE
      port map(D => \wsync1_rptr[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[14]_net_1\);
    
    \wbinaddr_RNI1ASQ2[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_3, S
         => \wbinaddr_RNI1ASQ2_S[4]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_4);
    
    \rgraynext[13]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIQTLC8_S[14]\, B => 
        \rbinaddr_RNI9QAU7_S[13]\, Y => \rgraynext[13]_net_1\);
    
    \wbinaddr[16]\ : SLE
      port map(D => \wbinaddr_2[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[16]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_57\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[17]_net_1\, B => 
        \rbinaddr_RNIJENN9_S[17]\, C => \rbinaddr_RNI8M26A_S[18]\, 
        D => fifo_empty_xhdl3_0_I_59_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[7]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[8]\);
    
    \rbinaddr_RNI14454[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_4, S
         => \rbinaddr_RNI14454_S[5]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_5);
    
    \rbinaddr[22]\ : SLE
      port map(D => \rbinaddr_3[22]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[22]_net_1\);
    
    \rddata_r_RNIQJIU[12]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[12]\, C => 
        \rddata_r[12]_net_1\, Y => N_283);
    
    \rsync1_wptr[1]\ : SLE
      port map(D => \waddr_gray[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[1]_net_1\);
    
    \rbinaddr_RNIV7C99[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_15, S
         => \rbinaddr_RNIV7C99_S[16]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_16);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_75\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[3]_net_1\, B => 
        \rbinaddr_RNI01753_S[3]\, C => \rbinaddr_RNI0I5L3_S[4]\, 
        D => fifo_empty_xhdl3_0_I_77_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[0]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[1]\);
    
    \rddata_r_RNIFC851[8]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[8]\, C => 
        \rddata_r[8]_net_1\, Y => N_435);
    
    \rgraynext[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI9QAU7_S[13]\, B => 
        \rbinaddr_RNIPNVF7_S[12]\, Y => \rgraynext[12]_net_1\);
    
    \raddr_gray[7]\ : SLE
      port map(D => \rgraynext[7]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[7]_net_1\);
    
    \wbinaddr_RNISS0M8[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_15, S
         => \wbinaddr_RNISS0M8_S[16]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_16);
    
    \rddata_r[1]\ : SLE
      port map(D => \port_xhdl7[1]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[1]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_99\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \rbinaddr_RNI79FFG_S[32]\, C
         => \rsync2_wptr[32]_net_1\, D => GND_net_1, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[15]\, S => OPEN, Y => OPEN, 
        FCO => fifo_empty_xhdl3_0_N_2);
    
    \waddr_gray[12]\ : SLE
      port map(D => \wgraynext[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[12]_net_1\);
    
    \rddata_r[6]\ : SLE
      port map(D => \port_xhdl7[6]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[6]_net_1\);
    
    \wbinaddr[9]\ : SLE
      port map(D => \wbinaddr_2[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[9]_net_1\);
    
    \rddata_r_RNI092O[60]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[60]\, C => 
        \rddata_r[60]_net_1\, Y => N_218);
    
    \rbinaddr_RNIA7F7E[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_26, S
         => \rbinaddr_RNIA7F7E_S[27]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_27);
    
    \wsync2_rptr[29]\ : SLE
      port map(D => \wsync1_rptr[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[29]_net_1\);
    
    \rsync1_wptr[29]\ : SLE
      port map(D => \waddr_gray[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[29]_net_1\);
    
    \rsync1_wptr[11]\ : SLE
      port map(D => \waddr_gray[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[11]_net_1\);
    
    \raddr_gray[4]\ : SLE
      port map(D => \rgraynext[4]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[4]_net_1\);
    
    \rddata_r[19]\ : SLE
      port map(D => \port_xhdl7[19]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[19]_net_1\);
    
    un13_writefull_0_I_93 : ARI1
      generic map(INIT => x"66900")

      port map(A => VCC_net_1, B => \wsync2_rptr[30]_net_1\, C
         => \wbinaddr_RNIUJD6A_S[31]\, D => 
        \wbinaddr_RNI9OB6A_S[30]\, FCI => 
        \un13_writefull_0_data_tmp[14]\, S => OPEN, Y => OPEN, 
        FCO => un13_writefull_0_N_2);
    
    \raddr_gray[30]\ : SLE
      port map(D => \rgraynext[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[30]_net_1\);
    
    \wsync2_rptr[19]\ : SLE
      port map(D => \wsync1_rptr[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[19]_net_1\);
    
    \rbinaddr_RNI79FFG[32]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[32]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_31, S
         => \rbinaddr_RNI79FFG_S[32]\, Y => OPEN, FCO => OPEN);
    
    \rddata_r_RNITMIU[15]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[15]\, C => 
        \rddata_r[15]_net_1\, Y => N_415);
    
    \rbinaddr_RNISAUDC[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_22, S
         => \rbinaddr_RNISAUDC_S[23]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_23);
    
    \rbinaddr[7]\ : SLE
      port map(D => \rbinaddr_3[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[7]_net_1\);
    
    \wbinaddr_RNIFP0M9[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_17, S
         => \wbinaddr_RNIFP0M9_S[18]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_18);
    
    un13_writefull_0_I_63 : ARI1
      generic map(INIT => x"60609")

      port map(A => \wsync2_rptr[21]_net_1\, B => 
        \wbinaddr_RNIHB26A_S[21]\, C => \wbinaddr_RNI6636A_S[22]\, 
        D => un13_writefull_0_N_27, FCI => 
        \un13_writefull_0_data_tmp[9]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[10]\);
    
    \rddata_r[16]\ : SLE
      port map(D => \port_xhdl7[16]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[16]_net_1\);
    
    \wsync2_rptr[23]\ : SLE
      port map(D => \wsync1_rptr[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[23]_net_1\);
    
    \waddr_gray[24]\ : SLE
      port map(D => \wgraynext[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[24]_net_1\);
    
    \rsync1_wptr[14]\ : SLE
      port map(D => \waddr_gray[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[14]_net_1\);
    
    \rddata_r_RNI85851[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[1]\, C => 
        \rddata_r[1]_net_1\, Y => N_150);
    
    \rddata_r[37]\ : SLE
      port map(D => \port_xhdl7[37]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[37]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[28]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI0HRLE_S[28]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[28]\);
    
    \rddata_r_RNIPIIU[11]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[11]\, C => 
        \rddata_r[11]_net_1\, Y => N_284);
    
    un13_writefull_0_I_81 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[27]_net_1\, B => 
        \wgraynext[26]_net_1\, C => \wgraynext[27]_net_1\, D => 
        \wsync2_rptr[26]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[12]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[13]\);
    
    \Read_Bin_Ptr.rbinaddr_3[0]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI6KBL1_S[0]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[0]\);
    
    \wsync2_rptr[13]\ : SLE
      port map(D => \wsync1_rptr[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[13]_net_1\);
    
    \rsync2_wptr[4]\ : SLE
      port map(D => \rsync1_wptr[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[4]_net_1\);
    
    \rsync2_wptr[16]\ : SLE
      port map(D => \rsync1_wptr[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[16]_net_1\);
    
    un13_writefull_0_I_1 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[1]_net_1\, B => 
        \wgraynext[0]_net_1\, C => \wgraynext[1]_net_1\, D => 
        \wsync2_rptr[0]_net_1\, FCI => GND_net_1, S => OPEN, Y
         => OPEN, FCO => \un13_writefull_0_data_tmp[0]\);
    
    \wgraynext[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIL3PD1_S[1]\, B => 
        \wbinaddr_RNIJ3OU_S[0]\, Y => \wgraynext[0]_net_1\);
    
    \wbinaddr_RNIN9167[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_12, S
         => \wbinaddr_RNIN9167_S[13]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_13);
    
    \rbinaddr[20]\ : SLE
      port map(D => \rbinaddr_3[20]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[20]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[30]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI9OB6A_S[30]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[30]\);
    
    \wsync1_rptr[5]\ : SLE
      port map(D => \raddr_gray[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[5]_net_1\);
    
    \wbinaddr_RNI2G1M6[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_11, S
         => \wbinaddr_RNI2G1M6_S[12]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_12);
    
    \rddata_r[57]\ : SLE
      port map(D => \port_xhdl7[57]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[57]_net_1\);
    
    \wsync2_rptr[21]\ : SLE
      port map(D => \wsync1_rptr[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[21]_net_1\);
    
    \rgraynext[31]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI79FFG_S[32]\, B => 
        \rbinaddr_RNIM321G_S[31]\, Y => \rgraynext[31]_net_1\);
    
    \rbinaddr[18]\ : SLE
      port map(D => \rbinaddr_3[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[18]_net_1\);
    
    fifo_empty_xhdl3_RNIA7D51 : ARI1
      generic map(INIT => x"400C4")

      port map(A => \fifo_empty_xhdl3\, B => N_98, C => 
        axi_current_state_0, D => N_72_i, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_rbinnext_cry_0_cy);
    
    \waddr_gray[0]\ : SLE
      port map(D => \wgraynext[0]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[0]_net_1\);
    
    \rsync1_wptr[9]\ : SLE
      port map(D => \waddr_gray[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[9]_net_1\);
    
    \rbinaddr_RNIQTLC8[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_13, S
         => \rbinaddr_RNIQTLC8_S[14]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_14);
    
    \wbinaddr_RNI9OB6A[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_29, S
         => \wbinaddr_RNI9OB6A_S[30]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_30);
    
    \wsync1_rptr[3]\ : SLE
      port map(D => \raddr_gray[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[3]_net_1\);
    
    \wsync2_rptr[11]\ : SLE
      port map(D => \wsync1_rptr[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[11]_net_1\);
    
    \rddata_r_RNI4C1O[55]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[55]\, C => 
        \rddata_r[55]_net_1\, Y => N_430);
    
    \wbinaddr_RNIHB26A[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_20, S
         => \wbinaddr_RNIHB26A_S[21]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_21);
    
    \Read_Bin_Ptr.rbinaddr_3[32]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI79FFG_S[32]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[32]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_93\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[5]_net_1\, B => 
        \rbinaddr_RNI14454_S[5]\, C => \rbinaddr_RNI3N2L4_S[6]\, 
        D => fifo_empty_xhdl3_0_I_95_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[1]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[2]\);
    
    \wbinaddr_RNIJU46A[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_23, S
         => \wbinaddr_RNIJU46A_S[24]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_24);
    
    \wsync1_rptr[32]\ : SLE
      port map(D => \raddr_gray[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[32]_net_1\);
    
    \wbinaddr_RNIUJD6A[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[31]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_30, S
         => \wbinaddr_RNIUJD6A_S[31]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_31);
    
    \rsync2_wptr[5]\ : SLE
      port map(D => \rsync1_wptr[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[5]_net_1\);
    
    \rbinaddr[12]\ : SLE
      port map(D => \rbinaddr_3[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[12]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[15]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI40168_S[15]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[15]\);
    
    \wsync1_rptr[31]\ : SLE
      port map(D => \raddr_gray[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[31]_net_1\);
    
    \rddata_r[27]\ : SLE
      port map(D => \port_xhdl7[27]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[27]_net_1\);
    
    \rddata_r_RNI3AVN[37]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[37]\, C => 
        \rddata_r[37]_net_1\, Y => N_426);
    
    \raddr_gray[22]\ : SLE
      port map(D => \rgraynext[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[22]_net_1\);
    
    \wsync1_rptr[7]\ : SLE
      port map(D => \raddr_gray[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[7]_net_1\);
    
    \wgraynext[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIEN166_S[11]\, B => 
        \wbinaddr_RNIRV1M5_S[10]\, Y => \wgraynext[10]_net_1\);
    
    \wbinaddr_RNIAP06A[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_18, S
         => \wbinaddr_RNIAP06A_S[19]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_19);
    
    un13_writefull_0_I_69 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[23]_net_1\, B => 
        \wgraynext[22]_net_1\, C => \wgraynext[23]_net_1\, D => 
        \wsync2_rptr[22]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[10]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[11]\);
    
    \rsync1_wptr[23]\ : SLE
      port map(D => \waddr_gray[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[23]_net_1\);
    
    \waddr_gray[15]\ : SLE
      port map(D => \wgraynext[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[15]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_71_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIB6IVB_S[22]\, B => 
        \rsync2_wptr[22]_net_1\, Y => fifo_empty_xhdl3_0_I_71_0);
    
    \wgraynext[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI1ASQ2_S[4]\, B => 
        \wbinaddr_RNIS6RB2_S[3]\, Y => \wgraynext[3]_net_1\);
    
    \rsync1_wptr[19]\ : SLE
      port map(D => \waddr_gray[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[19]_net_1\);
    
    \rddata_r[8]\ : SLE
      port map(D => \port_xhdl7[8]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[8]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[10]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIRV1M5_S[10]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[10]\);
    
    \rsync2_wptr[21]\ : SLE
      port map(D => \rsync1_wptr[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[21]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[1]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIL3PD1_S[1]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[1]\);
    
    \rddata_r_RNIU50O[41]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[41]\, C => 
        \rddata_r[41]_net_1\, Y => N_293);
    
    un13_writefull_0_I_21 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[7]_net_1\, B => 
        \wgraynext[6]_net_1\, C => \wgraynext[7]_net_1\, D => 
        \wsync2_rptr[6]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[2]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[3]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_51\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[11]_net_1\, B => 
        \rbinaddr_RNIAMK17_S[11]\, C => \rbinaddr_RNIPNVF7_S[12]\, 
        D => fifo_empty_xhdl3_0_I_53_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[5]\);
    
    fifo_empty_xhdl3 : SLE
      port map(D => fifo_empty_xhdl3_0_N_2_i, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_empty_xhdl3\);
    
    \raddr_gray[19]\ : SLE
      port map(D => \rgraynext[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[19]_net_1\);
    
    \raddr_gray[13]\ : SLE
      port map(D => \rgraynext[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[13]_net_1\);
    
    \wbinaddr_RNITH16A[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_19, S
         => \wbinaddr_RNITH16A_S[20]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_20);
    
    \rsync1_wptr[31]\ : SLE
      port map(D => \waddr_gray[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[31]_net_1\);
    
    \rgraynext[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI3N2L4_S[6]\, B => 
        \rbinaddr_RNI14454_S[5]\, Y => \rgraynext[5]_net_1\);
    
    \wbinaddr[7]\ : SLE
      port map(D => \wbinaddr_2[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[7]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[23]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIS146A_S[23]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[23]\);
    
    \waddr_gray[18]\ : SLE
      port map(D => \wgraynext[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[18]_net_1\);
    
    \rddata_r_RNI3TJU[29]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[29]\, C => 
        \rddata_r[29]_net_1\, Y => N_439);
    
    \wbinaddr_RNIO4QS1[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_1, S
         => \wbinaddr_RNIO4QS1_S[2]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_2);
    
    \wbinaddr[24]\ : SLE
      port map(D => \wbinaddr_2[24]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[24]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_17_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0HRLE_S[28]\, B => 
        \rsync2_wptr[28]_net_1\, Y => fifo_empty_xhdl3_0_I_17_0);
    
    \rbinaddr[3]\ : SLE
      port map(D => \rbinaddr_3[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[3]_net_1\);
    
    \raddr_gray[11]\ : SLE
      port map(D => \rgraynext[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[11]_net_1\);
    
    \rbinaddr[32]\ : SLE
      port map(D => \rbinaddr_3[32]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[32]_net_1\);
    
    \rbinaddr_RNIM321G[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[31]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_30, S
         => \rbinaddr_RNIM321G_S[31]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_31);
    
    \rbinaddr_RNILU2PD[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_25, S
         => \rbinaddr_RNILU2PD_S[26]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_26);
    
    \rddata_r[41]\ : SLE
      port map(D => \port_xhdl7[41]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[41]_net_1\);
    
    \rddata_r_RNI7F1O[58]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[58]\, C => 
        \rddata_r[58]_net_1\, Y => N_414);
    
    \wsync2_rptr[26]\ : SLE
      port map(D => \wsync1_rptr[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[26]_net_1\);
    
    \wgraynext[21]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI6636A_S[22]\, B => 
        \wbinaddr_RNIHB26A_S[21]\, Y => \wgraynext[21]_net_1\);
    
    \waddr_gray[27]\ : SLE
      port map(D => \wgraynext[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[27]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[29]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNINR74F_S[29]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[29]\);
    
    \rddata_r[40]\ : SLE
      port map(D => \port_xhdl7[40]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[40]_net_1\);
    
    \rbinaddr[10]\ : SLE
      port map(D => \rbinaddr_3[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[10]_net_1\);
    
    \waddr_gray[6]\ : SLE
      port map(D => \wgraynext[6]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[6]_net_1\);
    
    \wsync2_rptr[16]\ : SLE
      port map(D => \wsync1_rptr[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[16]_net_1\);
    
    \wgraynext[31]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIKGF6A_S[32]\, B => 
        \wbinaddr_RNIUJD6A_S[31]\, Y => \wgraynext[31]_net_1\);
    
    \rbinaddr_RNI6VKIF[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_29, S
         => \rbinaddr_RNI6VKIF_S[30]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_30);
    
    \rddata_r_RNIEB851[7]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[7]\, C => 
        \rddata_r[7]_net_1\, Y => N_434);
    
    \wsync2_rptr[5]\ : SLE
      port map(D => \wsync1_rptr[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[5]_net_1\);
    
    \wsync1_rptr[25]\ : SLE
      port map(D => \raddr_gray[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[25]_net_1\);
    
    \waddr_gray[3]\ : SLE
      port map(D => \wgraynext[3]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[3]_net_1\);
    
    \rbinaddr_RNI3N2L4[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_5, S
         => \rbinaddr_RNI3N2L4_S[6]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_6);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_59_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIV7C99_S[16]\, B => 
        \rsync2_wptr[16]_net_1\, Y => fifo_empty_xhdl3_0_I_59_0);
    
    \wgraynext[27]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIPR86A_S[28]\, B => 
        \wbinaddr_RNIUQ76A_S[27]\, Y => \wgraynext[27]_net_1\);
    
    \rddata_r_RNIT40O[40]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[40]\, C => 
        \rddata_r[40]_net_1\, Y => N_428);
    
    \wsync1_rptr[15]\ : SLE
      port map(D => \raddr_gray[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[15]_net_1\);
    
    \rsync2_wptr[24]\ : SLE
      port map(D => \rsync1_wptr[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[24]_net_1\);
    
    \rddata_r_RNI2RIU[19]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[19]\, C => 
        \rddata_r[19]_net_1\, Y => N_215);
    
    fifo_full_xhdl2 : SLE
      port map(D => \un9_writefull\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_full_xhdl2\);
    
    \wsync2_rptr[3]\ : SLE
      port map(D => \wsync1_rptr[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[3]_net_1\);
    
    \rbinaddr[2]\ : SLE
      port map(D => \rbinaddr_3[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[2]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[28]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIPR86A_S[28]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[28]\);
    
    \rsync1_wptr[8]\ : SLE
      port map(D => \waddr_gray[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[8]_net_1\);
    
    \rsync2_wptr[23]\ : SLE
      port map(D => \rsync1_wptr[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[23]_net_1\);
    
    \rsync2_wptr[7]\ : SLE
      port map(D => \rsync1_wptr[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[7]_net_1\);
    
    \rsync1_wptr[20]\ : SLE
      port map(D => \waddr_gray[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[20]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \waddr_gray[22]\ : SLE
      port map(D => \wgraynext[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[22]_net_1\);
    
    \rsync2_wptr[27]\ : SLE
      port map(D => \rsync1_wptr[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[27]_net_1\);
    
    \rgraynext[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIAMK17_S[11]\, B => 
        \rbinaddr_RNISL9J6_S[10]\, Y => \rgraynext[10]_net_1\);
    
    \rsync1_wptr[13]\ : SLE
      port map(D => \waddr_gray[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[13]_net_1\);
    
    \rbinaddr[6]\ : SLE
      port map(D => \rbinaddr_3[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[6]_net_1\);
    
    \rddata_r[17]\ : SLE
      port map(D => \port_xhdl7[17]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[17]_net_1\);
    
    \rbinaddr[30]\ : SLE
      port map(D => \rbinaddr_3[30]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[30]_net_1\);
    
    \wsync2_rptr[7]\ : SLE
      port map(D => \wsync1_rptr[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[7]_net_1\);
    
    \rddata_r[31]\ : SLE
      port map(D => \port_xhdl7[31]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[31]_net_1\);
    
    \rddata_r_RNI4C0O[47]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[47]\, C => 
        \rddata_r[47]_net_1\, Y => N_412);
    
    \rsync2_wptr[11]\ : SLE
      port map(D => \rsync1_wptr[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[11]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[12]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIPNVF7_S[12]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[12]\);
    
    \wsync1_rptr[27]\ : SLE
      port map(D => \raddr_gray[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[27]_net_1\);
    
    \raddr_gray[32]\ : SLE
      port map(D => \rbinaddr_RNI79FFG_S[32]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[32]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[4]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI0I5L3_S[4]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[4]\);
    
    \Read_Bin_Ptr.rbinaddr_3[30]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI6VKIF_S[30]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[30]\);
    
    \rddata_r[30]\ : SLE
      port map(D => \port_xhdl7[30]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[30]_net_1\);
    
    \rddata_r_RNI1QIU[18]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[18]\, C => 
        \rddata_r[18]_net_1\, Y => N_424);
    
    \rbinaddr_RNIEGASC[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_23, S
         => \rbinaddr_RNIEGASC_S[24]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_24);
    
    \wsync1_rptr[17]\ : SLE
      port map(D => \raddr_gray[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[17]_net_1\);
    
    \wbinaddr[3]\ : SLE
      port map(D => \wbinaddr_2[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[3]_net_1\);
    
    \rsync2_wptr[20]\ : SLE
      port map(D => \rsync1_wptr[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[20]_net_1\);
    
    \wgraynext[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIRV1M5_S[10]\, B => 
        \wbinaddr_RNI99265_S[9]\, Y => \wgraynext[9]_net_1\);
    
    \wsync1_rptr[30]\ : SLE
      port map(D => \raddr_gray[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[30]_net_1\);
    
    \wbinaddr[14]\ : SLE
      port map(D => \wbinaddr_2[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[14]_net_1\);
    
    \rsync1_wptr[6]\ : SLE
      port map(D => \waddr_gray[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[6]_net_1\);
    
    \wbinaddr_RNIBS56A[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_24, S
         => \wbinaddr_RNIBS56A_S[25]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_25);
    
    \Write_Bin_Ptr.wbinaddr_2[16]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNISS0M8_S[16]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[16]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_87\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[7]_net_1\, B => 
        \rbinaddr_RNI6B155_S[7]\, C => \rbinaddr_RNIA00L5_S[8]\, 
        D => fifo_empty_xhdl3_0_I_89_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[2]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[3]\);
    
    \raddr_gray[0]\ : SLE
      port map(D => \rgraynext[0]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[0]_net_1\);
    
    \rddata_r[51]\ : SLE
      port map(D => \port_xhdl7[51]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[51]_net_1\);
    
    \rddata_r_RNITMJU[23]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[23]\, C => 
        \rddata_r[23]_net_1\, Y => N_437);
    
    \rbinaddr_RNI1NMAD[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_24, S
         => \rbinaddr_RNI1NMAD_S[25]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_25);
    
    \waddr_gray[1]\ : SLE
      port map(D => \wgraynext[1]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[1]_net_1\);
    
    \rddata_r[50]\ : SLE
      port map(D => \port_xhdl7[50]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[50]_net_1\);
    
    \waddr_gray[5]\ : SLE
      port map(D => \wgraynext[5]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[5]_net_1\);
    
    \rbinaddr_RNI32A52[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_0, S
         => \rbinaddr_RNI32A52_S[1]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_1);
    
    \wbinaddr_RNIJ3OU[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_0_cy, 
        S => \wbinaddr_RNIJ3OU_S[0]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_0);
    
    \Read_Bin_Ptr.rbinaddr_3[17]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIJENN9_S[17]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[17]\);
    
    \wsync2_rptr[22]\ : SLE
      port map(D => \wsync1_rptr[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[22]_net_1\);
    
    \wsync2_rptr[30]\ : SLE
      port map(D => \wsync1_rptr[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[30]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[24]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIJU46A_S[24]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[24]\);
    
    \rbinaddr[29]\ : SLE
      port map(D => \rbinaddr_3[29]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[29]_net_1\);
    
    \rgraynext[21]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIB6IVB_S[22]\, B => 
        \rbinaddr_RNIR26HB_S[21]\, Y => \rgraynext[21]_net_1\);
    
    \rsync2_wptr[25]\ : SLE
      port map(D => \rsync1_wptr[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[25]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_53_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNISL9J6_S[10]\, B => 
        \rsync2_wptr[10]_net_1\, Y => fifo_empty_xhdl3_0_I_53_0);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_41_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIPNVF7_S[12]\, B => 
        \rsync2_wptr[12]_net_1\, Y => fifo_empty_xhdl3_0_I_41_0);
    
    \rgraynext[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNISL9J6_S[10]\, B => 
        \rbinaddr_RNIFMU46_S[9]\, Y => \rgraynext[9]_net_1\);
    
    \wsync2_rptr[12]\ : SLE
      port map(D => \wsync1_rptr[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[12]_net_1\);
    
    \rsync2_wptr[0]\ : SLE
      port map(D => \rsync1_wptr[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[0]_net_1\);
    
    \wsync1_rptr[4]\ : SLE
      port map(D => \raddr_gray[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[4]_net_1\);
    
    \wbinaddr[23]\ : SLE
      port map(D => \wbinaddr_2[23]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[23]_net_1\);
    
    \rddata_r[21]\ : SLE
      port map(D => \port_xhdl7[21]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[21]_net_1\);
    
    \rddata_r[0]\ : SLE
      port map(D => \port_xhdl7[0]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[0]_net_1\);
    
    \wgraynext[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIL3PD1_S[1]\, B => 
        \wbinaddr_RNIO4QS1_S[2]\, Y => \wgraynext[1]_net_1\);
    
    \wsync1_rptr[6]\ : SLE
      port map(D => \raddr_gray[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[6]_net_1\);
    
    \rgraynext[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI6B155_S[7]\, B => 
        \rbinaddr_RNI3N2L4_S[6]\, Y => \rgraynext[6]_net_1\);
    
    \wbinaddr[2]\ : SLE
      port map(D => \wbinaddr_2[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[2]_net_1\);
    
    \rsync1_wptr[26]\ : SLE
      port map(D => \waddr_gray[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[26]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[21]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIHB26A_S[21]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[21]\);
    
    \rddata_r[20]\ : SLE
      port map(D => \port_xhdl7[20]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[20]_net_1\);
    
    \rddata_r[4]\ : SLE
      port map(D => \port_xhdl7[4]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[4]_net_1\);
    
    \rsync2_wptr[14]\ : SLE
      port map(D => \rsync1_wptr[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[14]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[17]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNILQ069_S[17]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[17]\);
    
    \rsync2_wptr[13]\ : SLE
      port map(D => \rsync1_wptr[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[13]_net_1\);
    
    \wbinaddr_RNI7ET93[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_4, S
         => \wbinaddr_RNI7ET93_S[5]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_5);
    
    \wsync1_rptr[29]\ : SLE
      port map(D => \raddr_gray[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[29]_net_1\);
    
    \rbinaddr_RNI0I5L3[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_3, S
         => \rbinaddr_RNI0I5L3_S[4]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_4);
    
    \wbinaddr[6]\ : SLE
      port map(D => \wbinaddr_2[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[6]_net_1\);
    
    \rsync1_wptr[10]\ : SLE
      port map(D => \waddr_gray[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[10]_net_1\);
    
    \rgraynext[27]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0HRLE_S[28]\, B => 
        \rbinaddr_RNIA7F7E_S[27]\, Y => \rgraynext[27]_net_1\);
    
    \rsync2_wptr[17]\ : SLE
      port map(D => \rsync1_wptr[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[17]_net_1\);
    
    \rsync2_wptr[1]\ : SLE
      port map(D => \rsync1_wptr[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[1]_net_1\);
    
    \rddata_r_RNI2SJU[28]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[28]\, C => 
        \rddata_r[28]_net_1\, Y => N_210);
    
    \waddr_gray[25]\ : SLE
      port map(D => \wgraynext[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[25]_net_1\);
    
    \wsync1_rptr[19]\ : SLE
      port map(D => \raddr_gray[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[19]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[16]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIV7C99_S[16]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[16]\);
    
    \rddata_r[43]\ : SLE
      port map(D => \port_xhdl7[43]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[43]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_65_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIC0Q2B_S[20]\, B => 
        \rsync2_wptr[20]_net_1\, Y => fifo_empty_xhdl3_0_I_65_0);
    
    \wbinaddr_RNILQ069[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_16, S
         => \wbinaddr_RNILQ069_S[17]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_17);
    
    \Read_Bin_Ptr.rbinaddr_3[8]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIA00L5_S[8]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[8]\);
    
    \rddata_r_RNIUNJU[24]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[24]\, C => 
        \rddata_r[24]_net_1\, Y => N_425);
    
    \wsync2_rptr[25]\ : SLE
      port map(D => \wsync1_rptr[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[25]_net_1\);
    
    \rddata_r_RNI07VN[34]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[34]\, C => 
        \rddata_r[34]_net_1\, Y => N_158);
    
    \wgraynext[28]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNILT96A_S[29]\, B => 
        \wbinaddr_RNIPR86A_S[28]\, Y => \wgraynext[28]_net_1\);
    
    \rgraynext[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI01753_S[3]\, B => 
        \rbinaddr_RNI1H8L2_S[2]\, Y => \rgraynext[2]_net_1\);
    
    \waddr_gray[32]\ : SLE
      port map(D => \wbinaddr_RNIKGF6A_S[32]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[32]_net_1\);
    
    wren_2 : SLE
      port map(D => \wren_1\, CLK => SDRCLK_c, EN => 
        ahb_busyidle_cyc_i, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wren_2\);
    
    \raddr_gray[6]\ : SLE
      port map(D => \rgraynext[6]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[6]_net_1\);
    
    \raddr_gray[29]\ : SLE
      port map(D => \rgraynext[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[29]_net_1\);
    
    \raddr_gray[23]\ : SLE
      port map(D => \rgraynext[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[23]_net_1\);
    
    \wsync2_rptr[15]\ : SLE
      port map(D => \wsync1_rptr[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[15]_net_1\);
    
    \rsync2_wptr[31]\ : SLE
      port map(D => \rsync1_wptr[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[31]_net_1\);
    
    \rbinaddr_RNIR26HB[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_20, S
         => \rbinaddr_RNIR26HB_S[21]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_21);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_1\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[1]_net_1\, B => 
        \rbinaddr_RNI32A52_S[1]\, C => \rbinaddr_RNI1H8L2_S[2]\, 
        D => fifo_empty_xhdl3_0_I_5_0, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \fifo_empty_xhdl3_0_data_tmp[0]\);
    
    \Read_Bin_Ptr.rbinaddr_3[7]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI6B155_S[7]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[7]\);
    
    \waddr_gray[16]\ : SLE
      port map(D => \wgraynext[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[16]_net_1\);
    
    \waddr_gray[28]\ : SLE
      port map(D => \wgraynext[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[28]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[5]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI14454_S[5]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[5]\);
    
    \rsync2_wptr[10]\ : SLE
      port map(D => \rsync1_wptr[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[10]_net_1\);
    
    \wsync1_rptr[2]\ : SLE
      port map(D => \raddr_gray[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[2]_net_1\);
    
    \waddr_gray[2]\ : SLE
      port map(D => \wgraynext[2]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[2]_net_1\);
    
    un13_writefull_0_I_65 : CFG3
      generic map(INIT => x"96")

      port map(A => \wbinaddr_RNIHB26A_S[21]\, B => 
        \wsync2_rptr[20]_net_1\, C => \wbinaddr_RNITH16A_S[20]\, 
        Y => un13_writefull_0_N_27);
    
    \rddata_r[45]\ : SLE
      port map(D => \port_xhdl7[45]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[45]_net_1\);
    
    \raddr_gray[3]\ : SLE
      port map(D => \rgraynext[3]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[3]_net_1\);
    
    \raddr_gray[21]\ : SLE
      port map(D => \rgraynext[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[21]_net_1\);
    
    \wbinaddr_RNI6636A[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_21, S
         => \wbinaddr_RNI6636A_S[22]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_22);
    
    \rbinaddr[27]\ : SLE
      port map(D => \rbinaddr_3[27]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[27]_net_1\);
    
    \wsync1_rptr[0]\ : SLE
      port map(D => \raddr_gray[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[0]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[10]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNISL9J6_S[10]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[10]\);
    
    \rddata_r_RNISMKU[31]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[31]\, C => 
        \rddata_r[31]_net_1\, Y => N_209);
    
    \Read_Bin_Ptr.rbinaddr_3[6]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI3N2L4_S[6]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[6]\);
    
    \rbinaddr_RNI6KBL1[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_0_cy, 
        S => \rbinaddr_RNI6KBL1_S[0]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_0);
    
    rdinr_d : SLE
      port map(D => N_73_i_0, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdinr_d\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_95_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0I5L3_S[4]\, B => 
        \rsync2_wptr[4]_net_1\, Y => fifo_empty_xhdl3_0_I_95_0);
    
    \rgraynext[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI1H8L2_S[2]\, B => 
        \rbinaddr_RNI32A52_S[1]\, Y => \rgraynext[1]_net_1\);
    
    \rddata_r_RNIGD851[9]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[9]\, C => 
        \rddata_r[9]_net_1\, Y => N_286);
    
    \rbinaddr[4]\ : SLE
      port map(D => \rbinaddr_3[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[4]_net_1\);
    
    \rbinaddr_RNIPNVF7[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_11, S
         => \rbinaddr_RNIPNVF7_S[12]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_12);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_77_0\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI1H8L2_S[2]\, B => 
        \rsync2_wptr[2]_net_1\, Y => fifo_empty_xhdl3_0_I_77_0);
    
    \rddata_r_RNIA7851[3]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[3]\, C => 
        \rddata_r[3]_net_1\, Y => N_148);
    
    \Write_Bin_Ptr.wbinaddr_2[29]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNILT96A_S[29]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[29]\);
    
    \rsync1_wptr[3]\ : SLE
      port map(D => \waddr_gray[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[3]_net_1\);
    
    \rddata_r_RNI2A1O[53]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[53]\, C => 
        \rddata_r[53]_net_1\, Y => N_221);
    
    \Read_Bin_Ptr.rbinaddr_3[31]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIM321G_S[31]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[31]\);
    
    \rddata_r[48]\ : SLE
      port map(D => \port_xhdl7[48]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[48]_net_1\);
    
    \rbinaddr_RNIA00L5[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_7, S
         => \rbinaddr_RNIA00L5_S[8]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_8);
    
    \rddata_r_RNI6E1O[57]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[57]\, C => 
        \rddata_r[57]_net_1\, Y => N_413);
    
    \rddata_r_RNI3B1O[54]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[54]\, C => 
        \rddata_r[54]_net_1\, Y => N_429);
    
    \rddata_r[3]\ : SLE
      port map(D => \port_xhdl7[3]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[3]_net_1\);
    
    \rbinaddr[19]\ : SLE
      port map(D => \rbinaddr_3[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[19]_net_1\);
    
    \rsync2_wptr[15]\ : SLE
      port map(D => \rsync1_wptr[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[15]_net_1\);
    
    \wsync2_rptr[27]\ : SLE
      port map(D => \wsync1_rptr[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[27]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_81\ : ARI1
      generic map(INIT => x"62481")

      port map(A => \rsync2_wptr[9]_net_1\, B => 
        \rbinaddr_RNIFMU46_S[9]\, C => \rbinaddr_RNISL9J6_S[10]\, 
        D => fifo_empty_xhdl3_0_I_83_0, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[3]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[4]\);
    
    \wbinaddr[13]\ : SLE
      port map(D => \wbinaddr_2[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[13]_net_1\);
    
    \rddata_r_RNI3C2O[63]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[63]\, C => 
        \rddata_r[63]_net_1\, Y => N_217);
    
    \rddata_r[33]\ : SLE
      port map(D => \port_xhdl7[33]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[33]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[5]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI7ET93_S[5]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[5]\);
    
    \wsync2_rptr[4]\ : SLE
      port map(D => \wsync1_rptr[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[4]_net_1\);
    
    \rddata_r[11]\ : SLE
      port map(D => \port_xhdl7[11]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[11]_net_1\);
    
    \raddr_gray[15]\ : SLE
      port map(D => \rgraynext[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[15]_net_1\);
    
    \rsync1_wptr[16]\ : SLE
      port map(D => \waddr_gray[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[16]_net_1\);
    
    \wsync2_rptr[17]\ : SLE
      port map(D => \wsync1_rptr[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[17]_net_1\);
    
    \rddata_r_RNI4BVN[38]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[38]\, C => 
        \rddata_r[38]_net_1\, Y => N_410);
    
    \rddata_r_RNI190O[44]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[44]\, C => 
        \rddata_r[44]_net_1\, Y => N_290);
    
    \wsync2_rptr[6]\ : SLE
      port map(D => \wsync1_rptr[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[6]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[22]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIB6IVB_S[22]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[22]\);
    
    \rddata_r[10]\ : SLE
      port map(D => \port_xhdl7[10]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[10]_net_1\);
    
    \rddata_r[44]\ : SLE
      port map(D => \port_xhdl7[44]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[44]_net_1\);
    
    \rbinaddr_RNISL9J6[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_9, S
         => \rbinaddr_RNISL9J6_S[10]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_10);
    
    \rbinaddr_RNI9QAU7[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_12, S
         => \rbinaddr_RNI9QAU7_S[13]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_13);
    
    \raddr_gray[18]\ : SLE
      port map(D => \rgraynext[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[18]_net_1\);
    
    \rbinaddr_RNIC21R8[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_14, S
         => \rbinaddr_RNIC21R8_S[15]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_15);
    
    \wgraynext[26]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIUQ76A_S[27]\, B => 
        \wbinaddr_RNI4R66A_S[26]\, Y => \wgraynext[26]_net_1\);
    
    \wbinaddr[28]\ : SLE
      port map(D => \wbinaddr_2[28]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[28]_net_1\);
    
    \rsync2_wptr[9]\ : SLE
      port map(D => \rsync1_wptr[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[9]_net_1\);
    
    \rddata_r_RNIV61O[50]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[50]\, C => 
        \rddata_r[50]_net_1\, Y => N_420);
    
    \rddata_r[9]\ : SLE
      port map(D => \port_xhdl7[9]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[9]_net_1\);
    
    \wgraynext[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI2G1M6_S[12]\, B => 
        \wbinaddr_RNIEN166_S[11]\, Y => \wgraynext[11]_net_1\);
    
    \wbinaddr_RNIUQ76A[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_26, S
         => \wbinaddr_RNIUQ76A_S[27]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_27);
    
    \wbinaddr[29]\ : SLE
      port map(D => \wbinaddr_2[29]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[29]_net_1\);
    
    un9_writefull : CFG4
      generic map(INIT => x"0220")

      port map(A => \un7_writefull\, B => un13_writefull_0_N_2, C
         => \wsync2_rptr[32]_net_1\, D => 
        \wbinaddr_RNIKGF6A_S[32]\, Y => \un9_writefull\);
    
    \rddata_r[35]\ : SLE
      port map(D => \port_xhdl7[35]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[35]_net_1\);
    
    \rddata_r_RNIVOJU[25]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[25]\, C => 
        \rddata_r[25]_net_1\, Y => N_416);
    
    \rddata_r_RNISLIU[14]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[14]\, C => 
        \rddata_r[14]_net_1\, Y => N_281);
    
    \wsync2_rptr[31]\ : SLE
      port map(D => \wsync1_rptr[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[31]_net_1\);
    
    un13_writefull_0_I_87 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[29]_net_1\, B => 
        \wgraynext[28]_net_1\, C => \wgraynext[29]_net_1\, D => 
        \wsync2_rptr[28]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[13]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[14]\);
    
    \rsync1_wptr[22]\ : SLE
      port map(D => \waddr_gray[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[22]_net_1\);
    
    \rddata_r_RNIOHIU[10]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => \rdinr_d\, B => \port_xhdl7[10]\, C => 
        \rddata_r[10]_net_1\, Y => N_285);
    
    \wsync1_rptr[8]\ : SLE
      port map(D => \raddr_gray[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[8]_net_1\);
    
    \rsync2_wptr[22]\ : SLE
      port map(D => \rsync1_wptr[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[22]_net_1\);
    
    \rddata_r[53]\ : SLE
      port map(D => \port_xhdl7[53]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[53]_net_1\);
    
    \rsync1_wptr[30]\ : SLE
      port map(D => \waddr_gray[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[30]_net_1\);
    
    \rbinaddr_RNIUUDKA[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_18, S
         => \rbinaddr_RNIUUDKA_S[19]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_19);
    
    \Read_Bin_Ptr.rbinaddr_3[13]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI9QAU7_S[13]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[13]\);
    
    un13_writefull_0_I_33 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[11]_net_1\, B => 
        \wgraynext[10]_net_1\, C => \wgraynext[11]_net_1\, D => 
        \wsync2_rptr[10]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[4]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[5]\);
    
    \rbinaddr_RNI0HRLE[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_27, S
         => \rbinaddr_RNI0HRLE_S[28]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_28);
    
    \wbinaddr_RNID41M7[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_13, S
         => \wbinaddr_RNID41M7_S[14]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_14);
    
    \raddr_gray[1]\ : SLE
      port map(D => \rgraynext[1]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[1]_net_1\);
    
    \raddr_gray[5]\ : SLE
      port map(D => \rgraynext[5]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[5]_net_1\);
    
    \wbinaddr_RNIL3PD1[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un6_wbinnext_cry_0, S
         => \wbinaddr_RNIL3PD1_S[1]\, Y => OPEN, FCO => 
        un6_wbinnext_cry_1);
    
    \waddr_gray[19]\ : SLE
      port map(D => \wgraynext[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[19]_net_1\);
    
    \rddata_r[38]\ : SLE
      port map(D => \port_xhdl7[38]\, CLK => SDRCLK_c, EN => 
        \rdinr_d\, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rddata_r[38]_net_1\);
    
    \wgraynext[25]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI4R66A_S[26]\, B => 
        \wbinaddr_RNIBS56A_S[25]\, Y => \wgraynext[25]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_reset_syncHX_0 is

    port( SDRCLK_c  : in    std_logic;
          MSS_READY : in    std_logic;
          ARESET_n  : out   std_logic
        );

end CoreAHBLtoAXI_reset_syncHX_0;

architecture DEF_ARCH of CoreAHBLtoAXI_reset_syncHX_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \reset_sync_1\, \reset_sync_2\, VCC_net_1, GND_net_1
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    reset_sync_1_RNIGF7C : CLKINT
      port map(A => \reset_sync_1\, Y => ARESET_n);
    
    reset_sync_1 : SLE
      port map(D => \reset_sync_2\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => MSS_READY, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \reset_sync_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    reset_sync_2 : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => MSS_READY, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \reset_sync_2\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_rdch_ramHX is

    port( rdch_fifo_wr_data : in    std_logic_vector(31 downto 0);
          rdch_read_data    : out   std_logic_vector(31 downto 0);
          wbinaddr          : in    std_logic_vector(3 downto 0);
          rbinaddr          : in    std_logic_vector(3 downto 0);
          rdch_fifo_wr_en_r : in    std_logic;
          fifo_full_xhdl2   : in    std_logic;
          rdch_fifo_rd_en_r : in    std_logic;
          SDRCLK_c          : in    std_logic
        );

end CoreAHBLtoAXI_rdch_ramHX;

architecture DEF_ARCH of CoreAHBLtoAXI_rdch_ramHX is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component RAM64x18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_ADDR_CLK    : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ADDR_SRST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_ADDR_ARST_N : in    std_logic := 'U';
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_ADDR_EN     : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          B_ADDR_CLK    : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ADDR_SRST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_ADDR_ARST_N : in    std_logic := 'U';
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_ADDR_EN     : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_CLK         : in    std_logic := 'U';
          C_ADDR        : in    std_logic_vector(9 downto 0) := (others => 'U');
          C_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          C_WEN         : in    std_logic := 'U';
          C_BLK         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_ADDR_LAT    : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_EN          : in    std_logic := 'U';
          B_ADDR_LAT    : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          C_EN          : in    std_logic := 'U';
          C_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1, mem1_mem1_0_0_we, 
        mem1_mem1_0_1_we : std_logic;
    signal nc34, nc9, nc13, nc23, nc33, nc16, nc26, nc27, nc17, 
        nc36, nc37, nc5, nc4, nc25, nc15, nc35, nc28, nc18, nc38, 
        nc1, nc2, nc22, nc12, nc21, nc11, nc3, nc32, nc40, nc31, 
        nc7, nc6, nc19, nc29, nc39, nc8, nc20, nc10, nc24, nc14, 
        nc30 : std_logic;

begin 


    mem1_mem1_0_1_RNO : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_full_xhdl2, B => rdch_fifo_wr_en_r, Y
         => mem1_mem1_0_1_we);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    mem1_mem1_0_1 : RAM64x18
      port map(A_DOUT(17) => nc34, A_DOUT(16) => nc9, A_DOUT(15)
         => rdch_read_data(31), A_DOUT(14) => rdch_read_data(30), 
        A_DOUT(13) => rdch_read_data(29), A_DOUT(12) => 
        rdch_read_data(28), A_DOUT(11) => rdch_read_data(27), 
        A_DOUT(10) => rdch_read_data(26), A_DOUT(9) => 
        rdch_read_data(25), A_DOUT(8) => rdch_read_data(24), 
        A_DOUT(7) => rdch_read_data(23), A_DOUT(6) => 
        rdch_read_data(22), A_DOUT(5) => rdch_read_data(21), 
        A_DOUT(4) => rdch_read_data(20), A_DOUT(3) => 
        rdch_read_data(19), A_DOUT(2) => rdch_read_data(18), 
        A_DOUT(1) => rdch_read_data(17), A_DOUT(0) => 
        rdch_read_data(16), B_DOUT(17) => nc13, B_DOUT(16) => 
        nc23, B_DOUT(15) => nc33, B_DOUT(14) => nc16, B_DOUT(13)
         => nc26, B_DOUT(12) => nc27, B_DOUT(11) => nc17, 
        B_DOUT(10) => nc36, B_DOUT(9) => nc37, B_DOUT(8) => nc5, 
        B_DOUT(7) => nc4, B_DOUT(6) => nc25, B_DOUT(5) => nc15, 
        B_DOUT(4) => nc35, B_DOUT(3) => nc28, B_DOUT(2) => nc18, 
        B_DOUT(1) => nc38, B_DOUT(0) => nc1, BUSY => OPEN, 
        A_ADDR_CLK => VCC_net_1, A_DOUT_CLK => SDRCLK_c, 
        A_ADDR_SRST_N => VCC_net_1, A_DOUT_SRST_N => 
        rdch_fifo_rd_en_r, A_ADDR_ARST_N => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_ADDR_EN => VCC_net_1, 
        A_DOUT_EN => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_ADDR(9) => GND_net_1, A_ADDR(8) => 
        GND_net_1, A_ADDR(7) => rbinaddr(3), A_ADDR(6) => 
        rbinaddr(2), A_ADDR(5) => rbinaddr(1), A_ADDR(4) => 
        rbinaddr(0), A_ADDR(3) => GND_net_1, A_ADDR(2) => 
        GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, 
        B_ADDR_CLK => VCC_net_1, B_DOUT_CLK => SDRCLK_c, 
        B_ADDR_SRST_N => VCC_net_1, B_DOUT_SRST_N => 
        rdch_fifo_rd_en_r, B_ADDR_ARST_N => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_ADDR_EN => VCC_net_1, 
        B_DOUT_EN => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_ADDR(9) => GND_net_1, B_ADDR(8) => 
        GND_net_1, B_ADDR(7) => rbinaddr(3), B_ADDR(6) => 
        rbinaddr(2), B_ADDR(5) => rbinaddr(1), B_ADDR(4) => 
        rbinaddr(0), B_ADDR(3) => GND_net_1, B_ADDR(2) => 
        GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, 
        C_CLK => SDRCLK_c, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => wbinaddr(3), C_ADDR(6) => 
        wbinaddr(2), C_ADDR(5) => wbinaddr(1), C_ADDR(4) => 
        wbinaddr(0), C_ADDR(3) => GND_net_1, C_ADDR(2) => 
        GND_net_1, C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, 
        C_DIN(17) => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15)
         => rdch_fifo_wr_data(31), C_DIN(14) => 
        rdch_fifo_wr_data(30), C_DIN(13) => rdch_fifo_wr_data(29), 
        C_DIN(12) => rdch_fifo_wr_data(28), C_DIN(11) => 
        rdch_fifo_wr_data(27), C_DIN(10) => rdch_fifo_wr_data(26), 
        C_DIN(9) => rdch_fifo_wr_data(25), C_DIN(8) => 
        rdch_fifo_wr_data(24), C_DIN(7) => rdch_fifo_wr_data(23), 
        C_DIN(6) => rdch_fifo_wr_data(22), C_DIN(5) => 
        rdch_fifo_wr_data(21), C_DIN(4) => rdch_fifo_wr_data(20), 
        C_DIN(3) => rdch_fifo_wr_data(19), C_DIN(2) => 
        rdch_fifo_wr_data(18), C_DIN(1) => rdch_fifo_wr_data(17), 
        C_DIN(0) => rdch_fifo_wr_data(16), C_WEN => 
        mem1_mem1_0_1_we, C_BLK(1) => VCC_net_1, C_BLK(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_ADDR_LAT => VCC_net_1, 
        A_DOUT_LAT => GND_net_1, A_WIDTH(2) => VCC_net_1, 
        A_WIDTH(1) => GND_net_1, A_WIDTH(0) => GND_net_1, B_EN
         => GND_net_1, B_ADDR_LAT => VCC_net_1, B_DOUT_LAT => 
        GND_net_1, B_WIDTH(2) => VCC_net_1, B_WIDTH(1) => 
        GND_net_1, B_WIDTH(0) => GND_net_1, C_EN => VCC_net_1, 
        C_WIDTH(2) => VCC_net_1, C_WIDTH(1) => GND_net_1, 
        C_WIDTH(0) => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    mem1_mem1_0_0_RNO : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_full_xhdl2, B => rdch_fifo_wr_en_r, Y
         => mem1_mem1_0_0_we);
    
    mem1_mem1_0_0 : RAM64x18
      port map(A_DOUT(17) => nc2, A_DOUT(16) => nc22, A_DOUT(15)
         => rdch_read_data(15), A_DOUT(14) => rdch_read_data(14), 
        A_DOUT(13) => rdch_read_data(13), A_DOUT(12) => 
        rdch_read_data(12), A_DOUT(11) => rdch_read_data(11), 
        A_DOUT(10) => rdch_read_data(10), A_DOUT(9) => 
        rdch_read_data(9), A_DOUT(8) => rdch_read_data(8), 
        A_DOUT(7) => rdch_read_data(7), A_DOUT(6) => 
        rdch_read_data(6), A_DOUT(5) => rdch_read_data(5), 
        A_DOUT(4) => rdch_read_data(4), A_DOUT(3) => 
        rdch_read_data(3), A_DOUT(2) => rdch_read_data(2), 
        A_DOUT(1) => rdch_read_data(1), A_DOUT(0) => 
        rdch_read_data(0), B_DOUT(17) => nc12, B_DOUT(16) => nc21, 
        B_DOUT(15) => nc11, B_DOUT(14) => nc3, B_DOUT(13) => nc32, 
        B_DOUT(12) => nc40, B_DOUT(11) => nc31, B_DOUT(10) => nc7, 
        B_DOUT(9) => nc6, B_DOUT(8) => nc19, B_DOUT(7) => nc29, 
        B_DOUT(6) => nc39, B_DOUT(5) => nc8, B_DOUT(4) => nc20, 
        B_DOUT(3) => nc10, B_DOUT(2) => nc24, B_DOUT(1) => nc14, 
        B_DOUT(0) => nc30, BUSY => OPEN, A_ADDR_CLK => VCC_net_1, 
        A_DOUT_CLK => SDRCLK_c, A_ADDR_SRST_N => VCC_net_1, 
        A_DOUT_SRST_N => rdch_fifo_rd_en_r, A_ADDR_ARST_N => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_ADDR_EN => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(1) => VCC_net_1, 
        A_BLK(0) => VCC_net_1, A_ADDR(9) => GND_net_1, A_ADDR(8)
         => GND_net_1, A_ADDR(7) => rbinaddr(3), A_ADDR(6) => 
        rbinaddr(2), A_ADDR(5) => rbinaddr(1), A_ADDR(4) => 
        rbinaddr(0), A_ADDR(3) => GND_net_1, A_ADDR(2) => 
        GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, 
        B_ADDR_CLK => VCC_net_1, B_DOUT_CLK => SDRCLK_c, 
        B_ADDR_SRST_N => VCC_net_1, B_DOUT_SRST_N => 
        rdch_fifo_rd_en_r, B_ADDR_ARST_N => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_ADDR_EN => VCC_net_1, 
        B_DOUT_EN => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_ADDR(9) => GND_net_1, B_ADDR(8) => 
        GND_net_1, B_ADDR(7) => rbinaddr(3), B_ADDR(6) => 
        rbinaddr(2), B_ADDR(5) => rbinaddr(1), B_ADDR(4) => 
        rbinaddr(0), B_ADDR(3) => GND_net_1, B_ADDR(2) => 
        GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, 
        C_CLK => SDRCLK_c, C_ADDR(9) => GND_net_1, C_ADDR(8) => 
        GND_net_1, C_ADDR(7) => wbinaddr(3), C_ADDR(6) => 
        wbinaddr(2), C_ADDR(5) => wbinaddr(1), C_ADDR(4) => 
        wbinaddr(0), C_ADDR(3) => GND_net_1, C_ADDR(2) => 
        GND_net_1, C_ADDR(1) => GND_net_1, C_ADDR(0) => GND_net_1, 
        C_DIN(17) => GND_net_1, C_DIN(16) => GND_net_1, C_DIN(15)
         => rdch_fifo_wr_data(15), C_DIN(14) => 
        rdch_fifo_wr_data(14), C_DIN(13) => rdch_fifo_wr_data(13), 
        C_DIN(12) => rdch_fifo_wr_data(12), C_DIN(11) => 
        rdch_fifo_wr_data(11), C_DIN(10) => rdch_fifo_wr_data(10), 
        C_DIN(9) => rdch_fifo_wr_data(9), C_DIN(8) => 
        rdch_fifo_wr_data(8), C_DIN(7) => rdch_fifo_wr_data(7), 
        C_DIN(6) => rdch_fifo_wr_data(6), C_DIN(5) => 
        rdch_fifo_wr_data(5), C_DIN(4) => rdch_fifo_wr_data(4), 
        C_DIN(3) => rdch_fifo_wr_data(3), C_DIN(2) => 
        rdch_fifo_wr_data(2), C_DIN(1) => rdch_fifo_wr_data(1), 
        C_DIN(0) => rdch_fifo_wr_data(0), C_WEN => 
        mem1_mem1_0_0_we, C_BLK(1) => VCC_net_1, C_BLK(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_ADDR_LAT => VCC_net_1, 
        A_DOUT_LAT => GND_net_1, A_WIDTH(2) => VCC_net_1, 
        A_WIDTH(1) => GND_net_1, A_WIDTH(0) => GND_net_1, B_EN
         => GND_net_1, B_ADDR_LAT => VCC_net_1, B_DOUT_LAT => 
        GND_net_1, B_WIDTH(2) => VCC_net_1, B_WIDTH(1) => 
        GND_net_1, B_WIDTH(0) => GND_net_1, C_EN => VCC_net_1, 
        C_WIDTH(2) => VCC_net_1, C_WIDTH(1) => GND_net_1, 
        C_WIDTH(0) => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_RDCHANNELFIFOHX is

    port( rdch_read_data      : out   std_logic_vector(31 downto 0);
          rdch_fifo_wr_data   : in    std_logic_vector(31 downto 0);
          masterAddrInProg_0  : in    std_logic;
          valid_ahbcmd_i_o3_1 : in    std_logic;
          hsel2_0_a2_1        : in    std_logic;
          rdch_fifo_wr_en_r   : in    std_logic;
          rdch_fifo_rd_en_r   : in    std_logic;
          rdch_fifo_empty     : out   std_logic;
          SDRCLK_c            : in    std_logic;
          ARESET_n            : in    std_logic
        );

end CoreAHBLtoAXI_RDCHANNELFIFOHX;

architecture DEF_ARCH of CoreAHBLtoAXI_RDCHANNELFIFOHX is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CoreAHBLtoAXI_rdch_ramHX
    port( rdch_fifo_wr_data : in    std_logic_vector(31 downto 0) := (others => 'U');
          rdch_read_data    : out   std_logic_vector(31 downto 0);
          wbinaddr          : in    std_logic_vector(3 downto 0) := (others => 'U');
          rbinaddr          : in    std_logic_vector(3 downto 0) := (others => 'U');
          rdch_fifo_wr_en_r : in    std_logic := 'U';
          fifo_full_xhdl2   : in    std_logic := 'U';
          rdch_fifo_rd_en_r : in    std_logic := 'U';
          SDRCLK_c          : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal fifo_empty_xhdl3_0_N_2, fifo_empty_xhdl3_0_N_2_i, 
        \rbinaddr[18]_net_1\, VCC_net_1, \rbinaddr_3[18]\, 
        GND_net_1, \rbinaddr[19]_net_1\, \rbinaddr_3[19]\, 
        \rbinaddr[20]_net_1\, \rbinaddr_3[20]\, 
        \rbinaddr[21]_net_1\, \rbinaddr_3[21]\, 
        \rbinaddr[22]_net_1\, \rbinaddr_3[22]\, 
        \rbinaddr[23]_net_1\, \rbinaddr_3[23]\, 
        \rbinaddr[24]_net_1\, \rbinaddr_3[24]\, 
        \rbinaddr[25]_net_1\, \rbinaddr_3[25]\, 
        \rbinaddr[26]_net_1\, \rbinaddr_3[26]\, 
        \rbinaddr[27]_net_1\, \rbinaddr_3[27]\, 
        \rbinaddr[28]_net_1\, \rbinaddr_3[28]\, 
        \rbinaddr[29]_net_1\, \rbinaddr_3[29]\, 
        \rbinaddr[30]_net_1\, \rbinaddr_3[30]\, 
        \rbinaddr[31]_net_1\, \rbinaddr_3[31]\, 
        \rbinaddr[32]_net_1\, \rbinaddr_3[32]\, 
        \rbinaddr[3]_net_1\, \rbinaddr_3[3]\, \rbinaddr[4]_net_1\, 
        \rbinaddr_3[4]\, \rbinaddr[5]_net_1\, \rbinaddr_3[5]\, 
        \rbinaddr[6]_net_1\, \rbinaddr_3[6]\, \rbinaddr[7]_net_1\, 
        \rbinaddr_3[7]\, \rbinaddr[8]_net_1\, \rbinaddr_3[8]\, 
        \rbinaddr[9]_net_1\, \rbinaddr_3[9]\, 
        \rbinaddr[10]_net_1\, \rbinaddr_3[10]\, 
        \rbinaddr[11]_net_1\, \rbinaddr_3[11]\, 
        \rbinaddr[12]_net_1\, \rbinaddr_3[12]\, 
        \rbinaddr[13]_net_1\, \rbinaddr_3[13]\, 
        \rbinaddr[14]_net_1\, \rbinaddr_3[14]\, 
        \rbinaddr[15]_net_1\, \rbinaddr_3[15]\, 
        \rbinaddr[16]_net_1\, \rbinaddr_3[16]\, 
        \rbinaddr[17]_net_1\, \rbinaddr_3[17]\, 
        \rsync2_wptr[21]_net_1\, \rsync1_wptr[21]_net_1\, 
        \rsync2_wptr[22]_net_1\, \rsync1_wptr[22]_net_1\, 
        \rsync2_wptr[23]_net_1\, \rsync1_wptr[23]_net_1\, 
        \rsync2_wptr[24]_net_1\, \rsync1_wptr[24]_net_1\, 
        \rsync2_wptr[25]_net_1\, \rsync1_wptr[25]_net_1\, 
        \rsync2_wptr[26]_net_1\, \rsync1_wptr[26]_net_1\, 
        \rsync2_wptr[27]_net_1\, \rsync1_wptr[27]_net_1\, 
        \rsync2_wptr[28]_net_1\, \rsync1_wptr[28]_net_1\, 
        \rsync2_wptr[29]_net_1\, \rsync1_wptr[29]_net_1\, 
        \rsync2_wptr[30]_net_1\, \rsync1_wptr[30]_net_1\, 
        \rsync2_wptr[31]_net_1\, \rsync1_wptr[31]_net_1\, 
        \rsync2_wptr[32]_net_1\, \rsync1_wptr[32]_net_1\, 
        \rbinaddr[0]_net_1\, \rbinaddr_3[0]\, \rbinaddr[1]_net_1\, 
        \rbinaddr_3[1]\, \rbinaddr[2]_net_1\, \rbinaddr_3[2]\, 
        \rsync2_wptr[6]_net_1\, \rsync1_wptr[6]_net_1\, 
        \rsync2_wptr[7]_net_1\, \rsync1_wptr[7]_net_1\, 
        \rsync2_wptr[8]_net_1\, \rsync1_wptr[8]_net_1\, 
        \rsync2_wptr[9]_net_1\, \rsync1_wptr[9]_net_1\, 
        \rsync2_wptr[10]_net_1\, \rsync1_wptr[10]_net_1\, 
        \rsync2_wptr[11]_net_1\, \rsync1_wptr[11]_net_1\, 
        \rsync2_wptr[12]_net_1\, \rsync1_wptr[12]_net_1\, 
        \rsync2_wptr[13]_net_1\, \rsync1_wptr[13]_net_1\, 
        \rsync2_wptr[14]_net_1\, \rsync1_wptr[14]_net_1\, 
        \rsync2_wptr[15]_net_1\, \rsync1_wptr[15]_net_1\, 
        \rsync2_wptr[16]_net_1\, \rsync1_wptr[16]_net_1\, 
        \rsync2_wptr[17]_net_1\, \rsync1_wptr[17]_net_1\, 
        \rsync2_wptr[18]_net_1\, \rsync1_wptr[18]_net_1\, 
        \rsync2_wptr[19]_net_1\, \rsync1_wptr[19]_net_1\, 
        \rsync2_wptr[20]_net_1\, \rsync1_wptr[20]_net_1\, 
        \wsync2_rptr[24]_net_1\, \wsync1_rptr[24]_net_1\, 
        \wsync2_rptr[25]_net_1\, \wsync1_rptr[25]_net_1\, 
        \wsync2_rptr[26]_net_1\, \wsync1_rptr[26]_net_1\, 
        \wsync2_rptr[27]_net_1\, \wsync1_rptr[27]_net_1\, 
        \wsync2_rptr[28]_net_1\, \wsync1_rptr[28]_net_1\, 
        \wsync2_rptr[29]_net_1\, \wsync1_rptr[29]_net_1\, 
        \wsync2_rptr[30]_net_1\, \wsync1_rptr[30]_net_1\, 
        \wsync2_rptr[31]_net_1\, \wsync1_rptr[31]_net_1\, 
        \wsync2_rptr[32]_net_1\, \wsync1_rptr[32]_net_1\, 
        \rsync2_wptr[0]_net_1\, \rsync1_wptr[0]_net_1\, 
        \rsync2_wptr[1]_net_1\, \rsync1_wptr[1]_net_1\, 
        \rsync2_wptr[2]_net_1\, \rsync1_wptr[2]_net_1\, 
        \rsync2_wptr[3]_net_1\, \rsync1_wptr[3]_net_1\, 
        \rsync2_wptr[4]_net_1\, \rsync1_wptr[4]_net_1\, 
        \rsync2_wptr[5]_net_1\, \rsync1_wptr[5]_net_1\, 
        \wsync2_rptr[9]_net_1\, \wsync1_rptr[9]_net_1\, 
        \wsync2_rptr[10]_net_1\, \wsync1_rptr[10]_net_1\, 
        \wsync2_rptr[11]_net_1\, \wsync1_rptr[11]_net_1\, 
        \wsync2_rptr[12]_net_1\, \wsync1_rptr[12]_net_1\, 
        \wsync2_rptr[13]_net_1\, \wsync1_rptr[13]_net_1\, 
        \wsync2_rptr[14]_net_1\, \wsync1_rptr[14]_net_1\, 
        \wsync2_rptr[15]_net_1\, \wsync1_rptr[15]_net_1\, 
        \wsync2_rptr[16]_net_1\, \wsync1_rptr[16]_net_1\, 
        \wsync2_rptr[17]_net_1\, \wsync1_rptr[17]_net_1\, 
        \wsync2_rptr[18]_net_1\, \wsync1_rptr[18]_net_1\, 
        \wsync2_rptr[19]_net_1\, \wsync1_rptr[19]_net_1\, 
        \wsync2_rptr[20]_net_1\, \wsync1_rptr[20]_net_1\, 
        \wsync2_rptr[21]_net_1\, \wsync1_rptr[21]_net_1\, 
        \wsync2_rptr[22]_net_1\, \wsync1_rptr[22]_net_1\, 
        \wsync2_rptr[23]_net_1\, \wsync1_rptr[23]_net_1\, 
        \waddr_gray[27]_net_1\, \waddr_gray[28]_net_1\, 
        \waddr_gray[29]_net_1\, \waddr_gray[30]_net_1\, 
        \waddr_gray[31]_net_1\, \waddr_gray[32]_net_1\, 
        \wsync2_rptr[0]_net_1\, \wsync1_rptr[0]_net_1\, 
        \wsync2_rptr[1]_net_1\, \wsync1_rptr[1]_net_1\, 
        \wsync2_rptr[2]_net_1\, \wsync1_rptr[2]_net_1\, 
        \wsync2_rptr[3]_net_1\, \wsync1_rptr[3]_net_1\, 
        \wsync2_rptr[4]_net_1\, \wsync1_rptr[4]_net_1\, 
        \wsync2_rptr[5]_net_1\, \wsync1_rptr[5]_net_1\, 
        \wsync2_rptr[6]_net_1\, \wsync1_rptr[6]_net_1\, 
        \wsync2_rptr[7]_net_1\, \wsync1_rptr[7]_net_1\, 
        \wsync2_rptr[8]_net_1\, \wsync1_rptr[8]_net_1\, 
        \waddr_gray[12]_net_1\, \waddr_gray[13]_net_1\, 
        \waddr_gray[14]_net_1\, \waddr_gray[15]_net_1\, 
        \waddr_gray[16]_net_1\, \waddr_gray[17]_net_1\, 
        \waddr_gray[18]_net_1\, \waddr_gray[19]_net_1\, 
        \waddr_gray[20]_net_1\, \waddr_gray[21]_net_1\, 
        \waddr_gray[22]_net_1\, \waddr_gray[23]_net_1\, 
        \waddr_gray[24]_net_1\, \waddr_gray[25]_net_1\, 
        \waddr_gray[26]_net_1\, \raddr_gray[30]_net_1\, 
        \raddr_gray[31]_net_1\, \raddr_gray[32]_net_1\, 
        \waddr_gray[0]_net_1\, \waddr_gray[1]_net_1\, 
        \waddr_gray[2]_net_1\, \waddr_gray[3]_net_1\, 
        \waddr_gray[4]_net_1\, \waddr_gray[5]_net_1\, 
        \waddr_gray[6]_net_1\, \waddr_gray[7]_net_1\, 
        \waddr_gray[8]_net_1\, \waddr_gray[9]_net_1\, 
        \waddr_gray[10]_net_1\, \waddr_gray[11]_net_1\, 
        \raddr_gray[15]_net_1\, \raddr_gray[16]_net_1\, 
        \raddr_gray[17]_net_1\, \raddr_gray[18]_net_1\, 
        \raddr_gray[19]_net_1\, \raddr_gray[20]_net_1\, 
        \raddr_gray[21]_net_1\, \raddr_gray[22]_net_1\, 
        \raddr_gray[23]_net_1\, \raddr_gray[24]_net_1\, 
        \raddr_gray[25]_net_1\, \raddr_gray[26]_net_1\, 
        \raddr_gray[27]_net_1\, \raddr_gray[28]_net_1\, 
        \raddr_gray[29]_net_1\, \raddr_gray[0]_net_1\, 
        \raddr_gray[1]_net_1\, \raddr_gray[2]_net_1\, 
        \raddr_gray[3]_net_1\, \raddr_gray[4]_net_1\, 
        \raddr_gray[5]_net_1\, \raddr_gray[6]_net_1\, 
        \raddr_gray[7]_net_1\, \raddr_gray[8]_net_1\, 
        \raddr_gray[9]_net_1\, \raddr_gray[10]_net_1\, 
        \raddr_gray[11]_net_1\, \raddr_gray[12]_net_1\, 
        \raddr_gray[13]_net_1\, \raddr_gray[14]_net_1\, 
        \wgraynext[18]\, \wgraynext[19]\, \wgraynext[20]_net_1\, 
        \wgraynext[21]_net_1\, \wgraynext[22]_net_1\, 
        \wgraynext[23]_net_1\, \wgraynext[24]_net_1\, 
        \wgraynext[25]_net_1\, \wgraynext[26]_net_1\, 
        \wgraynext[27]_net_1\, \wgraynext[28]_net_1\, 
        \wgraynext[29]_net_1\, \wgraynext[30]_net_1\, 
        \wgraynext[31]_net_1\, \wbinaddr_RNIPD1S9_S[32]\, 
        \wgraynext[3]_net_1\, \wgraynext[4]_net_1\, 
        \wgraynext[5]_net_1\, \wgraynext[6]_net_1\, 
        \wgraynext[7]_net_1\, \wgraynext[8]_net_1\, 
        \wgraynext[9]_net_1\, \wgraynext[10]_net_1\, 
        \wgraynext[11]_net_1\, \wgraynext[12]_net_1\, 
        \wgraynext[13]_net_1\, \wgraynext[14]_net_1\, 
        \wgraynext[15]\, \wgraynext[16]\, \wgraynext[17]\, 
        \rgraynext[21]_net_1\, \rgraynext[22]_net_1\, 
        \rgraynext[23]_net_1\, \rgraynext[24]_net_1\, 
        \rgraynext[25]_net_1\, \rgraynext[26]_net_1\, 
        \rgraynext[27]_net_1\, \rgraynext[28]_net_1\, 
        \rgraynext[29]_net_1\, \rgraynext[30]_net_1\, 
        \rgraynext[31]_net_1\, \rbinaddr_RNIN7P39_S[32]\, 
        \wgraynext[0]_net_1\, \wgraynext[1]_net_1\, 
        \wgraynext[2]_net_1\, \rgraynext[6]_net_1\, 
        \rgraynext[7]_net_1\, \rgraynext[8]_net_1\, 
        \rgraynext[9]_net_1\, \rgraynext[10]_net_1\, 
        \rgraynext[11]_net_1\, \rgraynext[12]_net_1\, 
        \rgraynext[13]_net_1\, \rgraynext[14]_net_1\, 
        \rgraynext[15]_net_1\, \rgraynext[16]_net_1\, 
        \rgraynext[17]_net_1\, \rgraynext[18]_net_1\, 
        \rgraynext[19]_net_1\, \rgraynext[20]_net_1\, 
        \wbinaddr[24]_net_1\, \wbinaddr_2[24]\, 
        \wbinaddr[25]_net_1\, \wbinaddr_2[25]\, 
        \wbinaddr[26]_net_1\, \wbinaddr_2[26]\, 
        \wbinaddr[27]_net_1\, \wbinaddr_2[27]\, 
        \wbinaddr[28]_net_1\, \wbinaddr_2[28]\, 
        \wbinaddr[29]_net_1\, \wbinaddr_2[29]\, 
        \wbinaddr[30]_net_1\, \wbinaddr_2[30]\, 
        \wbinaddr[31]_net_1\, \wbinaddr_2[31]\, 
        \wbinaddr[32]_net_1\, \wbinaddr_2[32]\, 
        \rgraynext[0]_net_1\, \rgraynext[1]_net_1\, 
        \rgraynext[2]_net_1\, \rgraynext[3]_net_1\, 
        \rgraynext[4]_net_1\, \rgraynext[5]_net_1\, 
        \wbinaddr[9]_net_1\, \wbinaddr_2[9]\, 
        \wbinaddr[10]_net_1\, \wbinaddr_2[10]\, 
        \wbinaddr[11]_net_1\, \wbinaddr_2[11]\, 
        \wbinaddr[12]_net_1\, \wbinaddr_2[12]\, 
        \wbinaddr[13]_net_1\, \wbinaddr_2[13]\, 
        \wbinaddr[14]_net_1\, \wbinaddr_2[14]\, 
        \wbinaddr[15]_net_1\, \wbinaddr_2[15]\, 
        \wbinaddr[16]_net_1\, \wbinaddr_2[16]\, 
        \wbinaddr[17]_net_1\, \wbinaddr_2[17]\, 
        \wbinaddr[18]_net_1\, \wbinaddr_2[18]\, 
        \wbinaddr[19]_net_1\, \wbinaddr_2[19]\, 
        \wbinaddr[20]_net_1\, \wbinaddr_2[20]\, 
        \wbinaddr[21]_net_1\, \wbinaddr_2[21]\, 
        \wbinaddr[22]_net_1\, \wbinaddr_2[22]\, 
        \wbinaddr[23]_net_1\, \wbinaddr_2[23]\, 
        \wbinaddr[0]_net_1\, \wbinaddr_2[0]\, \wbinaddr[1]_net_1\, 
        \wbinaddr_2[1]\, \wbinaddr[2]_net_1\, \wbinaddr_2[2]\, 
        \wbinaddr[3]_net_1\, \wbinaddr_2[3]\, \wbinaddr[4]_net_1\, 
        \wbinaddr_2[4]\, \wbinaddr[5]_net_1\, \wbinaddr_2[5]\, 
        \wbinaddr[6]_net_1\, \wbinaddr_2[6]\, \wbinaddr[7]_net_1\, 
        \wbinaddr_2[7]\, \wbinaddr[8]_net_1\, \wbinaddr_2[8]\, 
        \rdch_fifo_empty\, \fifo_full_xhdl2\, un9_writefull_0, 
        un3_rbinnext_cry_0_cy, un3_rbinnext_cry_0, 
        \rbinaddr_RNIMQJL_S[0]\, un3_rbinnext_cry_1, 
        \rbinaddr_RNI0EAP_S[1]\, un3_rbinnext_cry_2, 
        \rbinaddr_RNIB21T_S[2]\, un3_rbinnext_cry_3, 
        \rbinaddr_RNINNN01_S[3]\, un3_rbinnext_cry_4, 
        \rbinaddr_RNI4EE41_S[4]\, un3_rbinnext_cry_5, 
        \rbinaddr_RNII5581_S[5]\, un3_rbinnext_cry_6, 
        \rbinaddr_RNI1URB1_S[6]\, un3_rbinnext_cry_7, 
        \rbinaddr_RNIHNIF1_S[7]\, un3_rbinnext_cry_8, 
        \rbinaddr_RNI2I9J1_S[8]\, un3_rbinnext_cry_9, 
        \rbinaddr_RNIKD0N1_S[9]\, un3_rbinnext_cry_10, 
        \rbinaddr_RNIEV812_S[10]\, un3_rbinnext_cry_11, 
        \rbinaddr_RNI9IHB2_S[11]\, un3_rbinnext_cry_12, 
        \rbinaddr_RNI56QL2_S[12]\, un3_rbinnext_cry_13, 
        \rbinaddr_RNI2R203_S[13]\, un3_rbinnext_cry_14, 
        \rbinaddr_RNI0HBA3_S[14]\, un3_rbinnext_cry_15, 
        \rbinaddr_RNIV7KK3_S[15]\, un3_rbinnext_cry_16, 
        \rbinaddr_RNIVVSU3_S[16]\, un3_rbinnext_cry_17, 
        \rbinaddr_RNI0P594_S[17]\, un3_rbinnext_cry_18, 
        \rbinaddr_RNI2JEJ4_S[18]\, un3_rbinnext_cry_19, 
        \rbinaddr_RNI5ENT4_S[19]\, un3_rbinnext_cry_20, 
        \rbinaddr_RNI02185_S[20]\, un3_rbinnext_cry_21, 
        \rbinaddr_RNISMAI5_S[21]\, un3_rbinnext_cry_22, 
        \rbinaddr_RNIPCKS5_S[22]\, un3_rbinnext_cry_23, 
        \rbinaddr_RNIN3U66_S[23]\, un3_rbinnext_cry_24, 
        \rbinaddr_RNIMR7H6_S[24]\, un3_rbinnext_cry_25, 
        \rbinaddr_RNIMKHR6_S[25]\, un3_rbinnext_cry_26, 
        \rbinaddr_RNINER57_S[26]\, un3_rbinnext_cry_27, 
        \rbinaddr_RNIP95G7_S[27]\, un3_rbinnext_cry_28, 
        \rbinaddr_RNIS5FQ7_S[28]\, un3_rbinnext_cry_29, 
        \rbinaddr_RNI03P48_S[29]\, un3_rbinnext_cry_30, 
        \rbinaddr_RNISO3F8_S[30]\, un3_rbinnext_cry_31, 
        \rbinaddr_RNIPFEP8_S[31]\, un3_wbinnext_cry_0_cy, 
        un3_wbinnext_cry_0, \wbinaddr_RNIO88G_S[0]\, 
        un3_wbinnext_cry_1, \wbinaddr_RNI7E1J_S[1]\, 
        un3_wbinnext_cry_2, \wbinaddr_RNINKQL_S[2]\, 
        un3_wbinnext_cry_3, \wbinaddr_RNI8SJO_S[3]\, 
        un3_wbinnext_cry_4, \wbinaddr_RNIQ4DR_S[4]\, 
        un3_wbinnext_cry_5, \wbinaddr_RNIDE6U_S[5]\, 
        un3_wbinnext_cry_6, \wbinaddr_RNI1PV01_S[6]\, 
        un3_wbinnext_cry_7, \wbinaddr_RNIM4P31_S[7]\, 
        un3_wbinnext_cry_8, \wbinaddr_RNICHI61_S[8]\, 
        un3_wbinnext_cry_9, \wbinaddr_RNI3VB91_S[9]\, 
        un3_wbinnext_cry_10, \wbinaddr_RNI289L1_S[10]\, 
        un3_wbinnext_cry_11, \wbinaddr_RNI2I612_S[11]\, 
        un3_wbinnext_cry_12, \wbinaddr_RNI3T3D2_S[12]\, 
        un3_wbinnext_cry_13, \wbinaddr_RNI591P2_S[13]\, 
        un3_wbinnext_cry_14, \wbinaddr_RNI8MU43_S[14]\, 
        un3_wbinnext_cry_15, \wbinaddr_RNIC4SG3_S[15]\, 
        un3_wbinnext_cry_16, \wbinaddr_RNIHJPS3_S[16]\, 
        un3_wbinnext_cry_17, \wbinaddr_RNIN3N84_S[17]\, 
        un3_wbinnext_cry_18, \wbinaddr_RNIUKKK4_S[18]\, 
        un3_wbinnext_cry_19, \wbinaddr_RNI67I05_S[19]\, 
        un3_wbinnext_cry_20, \wbinaddr_RNI6IGC5_S[20]\, 
        un3_wbinnext_cry_21, \wbinaddr_RNI7UEO5_S[21]\, 
        un3_wbinnext_cry_22, \wbinaddr_RNI9BD46_S[22]\, 
        un3_wbinnext_cry_23, \wbinaddr_RNICPBG6_S[23]\, 
        un3_wbinnext_cry_24, \wbinaddr_RNIG8AS6_S[24]\, 
        un3_wbinnext_cry_25, \wbinaddr_RNILO887_S[25]\, 
        un3_wbinnext_cry_26, \wbinaddr_RNIR97K7_S[26]\, 
        un3_wbinnext_cry_27, \wbinaddr_RNI2S508_S[27]\, 
        un3_wbinnext_cry_28, \wbinaddr_RNIAF4C8_S[28]\, 
        un3_wbinnext_cry_29, \wbinaddr_RNIJ33O8_S[29]\, 
        un3_wbinnext_cry_30, \wbinaddr_RNIKG249_S[30]\, 
        un3_wbinnext_cry_31, \wbinaddr_RNIMU1G9_S[31]\, 
        \fifo_empty_xhdl3_0_data_tmp[0]\, fifo_empty_xhdl3_0_N_81, 
        \fifo_empty_xhdl3_0_data_tmp[1]\, fifo_empty_xhdl3_0_N_21, 
        \fifo_empty_xhdl3_0_data_tmp[2]\, fifo_empty_xhdl3_0_N_6, 
        \fifo_empty_xhdl3_0_data_tmp[3]\, fifo_empty_xhdl3_0_N_11, 
        \fifo_empty_xhdl3_0_data_tmp[4]\, fifo_empty_xhdl3_0_N_16, 
        \fifo_empty_xhdl3_0_data_tmp[5]\, fifo_empty_xhdl3_0_N_41, 
        \fifo_empty_xhdl3_0_data_tmp[6]\, fifo_empty_xhdl3_0_N_51, 
        \fifo_empty_xhdl3_0_data_tmp[7]\, fifo_empty_xhdl3_0_N_46, 
        \fifo_empty_xhdl3_0_data_tmp[8]\, fifo_empty_xhdl3_0_N_36, 
        \fifo_empty_xhdl3_0_data_tmp[9]\, fifo_empty_xhdl3_0_N_61, 
        \fifo_empty_xhdl3_0_data_tmp[10]\, 
        fifo_empty_xhdl3_0_N_31, 
        \fifo_empty_xhdl3_0_data_tmp[11]\, 
        fifo_empty_xhdl3_0_N_26, 
        \fifo_empty_xhdl3_0_data_tmp[12]\, 
        fifo_empty_xhdl3_0_N_56, 
        \fifo_empty_xhdl3_0_data_tmp[13]\, 
        fifo_empty_xhdl3_0_N_66, 
        \fifo_empty_xhdl3_0_data_tmp[14]\, 
        fifo_empty_xhdl3_0_N_71, 
        \fifo_empty_xhdl3_0_data_tmp[15]\, 
        fifo_empty_xhdl3_0_N_76, \un13_writefull_0_data_tmp[0]\, 
        \un13_writefull_0_data_tmp[1]\, 
        \un13_writefull_0_data_tmp[2]\, 
        \un13_writefull_0_data_tmp[3]\, 
        \un13_writefull_0_data_tmp[4]\, 
        \un13_writefull_0_data_tmp[5]\, 
        \un13_writefull_0_data_tmp[6]\, 
        \un13_writefull_0_data_tmp[7]\, 
        \un13_writefull_0_data_tmp[8]\, 
        \un13_writefull_0_data_tmp[9]\, 
        \un13_writefull_0_data_tmp[10]\, 
        \un13_writefull_0_data_tmp[11]\, 
        \un13_writefull_0_data_tmp[12]\, 
        \un13_writefull_0_data_tmp[13]\, 
        \un13_writefull_0_data_tmp[14]\, un13_writefull_0_N_2, 
        \un7_writefull\ : std_logic;

    for all : CoreAHBLtoAXI_rdch_ramHX
	Use entity work.CoreAHBLtoAXI_rdch_ramHX(DEF_ARCH);
begin 

    rdch_fifo_empty <= \rdch_fifo_empty\;

    \waddr_gray[31]\ : SLE
      port map(D => \wgraynext[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[31]_net_1\);
    
    \rbinaddr_RNI56QL2[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_11, S
         => \rbinaddr_RNI56QL2_S[12]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_12);
    
    \rbinaddr_RNI5ENT4[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_18, S
         => \rbinaddr_RNI5ENT4_S[19]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_19);
    
    \rbinaddr[29]\ : SLE
      port map(D => \rbinaddr_3[29]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[29]_net_1\);
    
    \rsync2_wptr[19]\ : SLE
      port map(D => \rsync1_wptr[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[19]_net_1\);
    
    \raddr_gray[25]\ : SLE
      port map(D => \rgraynext[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[25]_net_1\);
    
    \rbinaddr[14]\ : SLE
      port map(D => \rbinaddr_3[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[14]_net_1\);
    
    \rbinaddr_RNIMQJL[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_0_cy, 
        S => \rbinaddr_RNIMQJL_S[0]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_0);
    
    \wbinaddr[31]\ : SLE
      port map(D => \wbinaddr_2[31]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[31]_net_1\);
    
    \waddr_gray[14]\ : SLE
      port map(D => \wgraynext[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[14]_net_1\);
    
    \rsync1_wptr[30]\ : SLE
      port map(D => \waddr_gray[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[30]_net_1\);
    
    \rbinaddr[27]\ : SLE
      port map(D => \rbinaddr_3[27]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[27]_net_1\);
    
    \waddr_gray[22]\ : SLE
      port map(D => \wgraynext[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[22]_net_1\);
    
    \rsync2_wptr[32]\ : SLE
      port map(D => \rsync1_wptr[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[32]_net_1\);
    
    \wbinaddr_RNIAF4C8[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_27, S
         => \wbinaddr_RNIAF4C8_S[28]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_28);
    
    \rsync2_wptr[15]\ : SLE
      port map(D => \rsync1_wptr[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[15]_net_1\);
    
    \wsync1_rptr[27]\ : SLE
      port map(D => \raddr_gray[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[27]_net_1\);
    
    \wbinaddr[13]\ : SLE
      port map(D => \wbinaddr_2[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[13]_net_1\);
    
    \raddr_gray[0]\ : SLE
      port map(D => \rgraynext[0]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[0]_net_1\);
    
    \wbinaddr_RNIDE6U[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_4, S
         => \wbinaddr_RNIDE6U_S[5]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_5);
    
    \raddr_gray[3]\ : SLE
      port map(D => \rgraynext[3]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[3]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_21\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[26]_net_1\, B => 
        \rbinaddr_RNINER57_S[26]\, C => \rbinaddr_RNIP95G7_S[27]\, 
        D => fifo_empty_xhdl3_0_N_66, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[12]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[13]\);
    
    \rgraynext[14]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIV7KK3_S[15]\, B => 
        \rbinaddr_RNI0HBA3_S[14]\, Y => \rgraynext[14]_net_1\);
    
    \rsync2_wptr[8]\ : SLE
      port map(D => \rsync1_wptr[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[8]_net_1\);
    
    \wbinaddr[3]\ : SLE
      port map(D => \wbinaddr_2[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[3]_net_1\);
    
    U_RDCH_RAM : CoreAHBLtoAXI_rdch_ramHX
      port map(rdch_fifo_wr_data(31) => rdch_fifo_wr_data(31), 
        rdch_fifo_wr_data(30) => rdch_fifo_wr_data(30), 
        rdch_fifo_wr_data(29) => rdch_fifo_wr_data(29), 
        rdch_fifo_wr_data(28) => rdch_fifo_wr_data(28), 
        rdch_fifo_wr_data(27) => rdch_fifo_wr_data(27), 
        rdch_fifo_wr_data(26) => rdch_fifo_wr_data(26), 
        rdch_fifo_wr_data(25) => rdch_fifo_wr_data(25), 
        rdch_fifo_wr_data(24) => rdch_fifo_wr_data(24), 
        rdch_fifo_wr_data(23) => rdch_fifo_wr_data(23), 
        rdch_fifo_wr_data(22) => rdch_fifo_wr_data(22), 
        rdch_fifo_wr_data(21) => rdch_fifo_wr_data(21), 
        rdch_fifo_wr_data(20) => rdch_fifo_wr_data(20), 
        rdch_fifo_wr_data(19) => rdch_fifo_wr_data(19), 
        rdch_fifo_wr_data(18) => rdch_fifo_wr_data(18), 
        rdch_fifo_wr_data(17) => rdch_fifo_wr_data(17), 
        rdch_fifo_wr_data(16) => rdch_fifo_wr_data(16), 
        rdch_fifo_wr_data(15) => rdch_fifo_wr_data(15), 
        rdch_fifo_wr_data(14) => rdch_fifo_wr_data(14), 
        rdch_fifo_wr_data(13) => rdch_fifo_wr_data(13), 
        rdch_fifo_wr_data(12) => rdch_fifo_wr_data(12), 
        rdch_fifo_wr_data(11) => rdch_fifo_wr_data(11), 
        rdch_fifo_wr_data(10) => rdch_fifo_wr_data(10), 
        rdch_fifo_wr_data(9) => rdch_fifo_wr_data(9), 
        rdch_fifo_wr_data(8) => rdch_fifo_wr_data(8), 
        rdch_fifo_wr_data(7) => rdch_fifo_wr_data(7), 
        rdch_fifo_wr_data(6) => rdch_fifo_wr_data(6), 
        rdch_fifo_wr_data(5) => rdch_fifo_wr_data(5), 
        rdch_fifo_wr_data(4) => rdch_fifo_wr_data(4), 
        rdch_fifo_wr_data(3) => rdch_fifo_wr_data(3), 
        rdch_fifo_wr_data(2) => rdch_fifo_wr_data(2), 
        rdch_fifo_wr_data(1) => rdch_fifo_wr_data(1), 
        rdch_fifo_wr_data(0) => rdch_fifo_wr_data(0), 
        rdch_read_data(31) => rdch_read_data(31), 
        rdch_read_data(30) => rdch_read_data(30), 
        rdch_read_data(29) => rdch_read_data(29), 
        rdch_read_data(28) => rdch_read_data(28), 
        rdch_read_data(27) => rdch_read_data(27), 
        rdch_read_data(26) => rdch_read_data(26), 
        rdch_read_data(25) => rdch_read_data(25), 
        rdch_read_data(24) => rdch_read_data(24), 
        rdch_read_data(23) => rdch_read_data(23), 
        rdch_read_data(22) => rdch_read_data(22), 
        rdch_read_data(21) => rdch_read_data(21), 
        rdch_read_data(20) => rdch_read_data(20), 
        rdch_read_data(19) => rdch_read_data(19), 
        rdch_read_data(18) => rdch_read_data(18), 
        rdch_read_data(17) => rdch_read_data(17), 
        rdch_read_data(16) => rdch_read_data(16), 
        rdch_read_data(15) => rdch_read_data(15), 
        rdch_read_data(14) => rdch_read_data(14), 
        rdch_read_data(13) => rdch_read_data(13), 
        rdch_read_data(12) => rdch_read_data(12), 
        rdch_read_data(11) => rdch_read_data(11), 
        rdch_read_data(10) => rdch_read_data(10), 
        rdch_read_data(9) => rdch_read_data(9), rdch_read_data(8)
         => rdch_read_data(8), rdch_read_data(7) => 
        rdch_read_data(7), rdch_read_data(6) => rdch_read_data(6), 
        rdch_read_data(5) => rdch_read_data(5), rdch_read_data(4)
         => rdch_read_data(4), rdch_read_data(3) => 
        rdch_read_data(3), rdch_read_data(2) => rdch_read_data(2), 
        rdch_read_data(1) => rdch_read_data(1), rdch_read_data(0)
         => rdch_read_data(0), wbinaddr(3) => \wbinaddr[3]_net_1\, 
        wbinaddr(2) => \wbinaddr[2]_net_1\, wbinaddr(1) => 
        \wbinaddr[1]_net_1\, wbinaddr(0) => \wbinaddr[0]_net_1\, 
        rbinaddr(3) => \rbinaddr[3]_net_1\, rbinaddr(2) => 
        \rbinaddr[2]_net_1\, rbinaddr(1) => \rbinaddr[1]_net_1\, 
        rbinaddr(0) => \rbinaddr[0]_net_1\, rdch_fifo_wr_en_r => 
        rdch_fifo_wr_en_r, fifo_full_xhdl2 => \fifo_full_xhdl2\, 
        rdch_fifo_rd_en_r => rdch_fifo_rd_en_r, SDRCLK_c => 
        SDRCLK_c);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_52\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI56QL2_S[12]\, B => 
        \rsync2_wptr[11]_net_1\, C => \rbinaddr_RNI9IHB2_S[11]\, 
        Y => fifo_empty_xhdl3_0_N_41);
    
    \Write_Bin_Ptr.wbinaddr_2[28]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIAF4C8_S[28]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[28]\);
    
    \wbinaddr[28]\ : SLE
      port map(D => \wbinaddr_2[28]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[28]_net_1\);
    
    \rsync2_wptr[28]\ : SLE
      port map(D => \rsync1_wptr[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[28]_net_1\);
    
    \wgraynext[25]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIR97K7_S[26]\, B => 
        \wbinaddr_RNILO887_S[25]\, Y => \wgraynext[25]_net_1\);
    
    \wbinaddr[9]\ : SLE
      port map(D => \wbinaddr_2[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[9]_net_1\);
    
    un13_writefull_0_I_93 : ARI1
      generic map(INIT => x"66900")

      port map(A => VCC_net_1, B => \wsync2_rptr[30]_net_1\, C
         => \wbinaddr_RNIMU1G9_S[31]\, D => 
        \wbinaddr_RNIKG249_S[30]\, FCI => 
        \un13_writefull_0_data_tmp[14]\, S => OPEN, Y => OPEN, 
        FCO => un13_writefull_0_N_2);
    
    \wgraynext[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI3VB91_S[9]\, B => 
        \wbinaddr_RNICHI61_S[8]\, Y => \wgraynext[8]_net_1\);
    
    \rbinaddr[32]\ : SLE
      port map(D => \rbinaddr_3[32]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[32]_net_1\);
    
    \wgraynext[20]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI7UEO5_S[21]\, B => 
        \wbinaddr_RNI6IGC5_S[20]\, Y => \wgraynext[20]_net_1\);
    
    \rsync1_wptr[15]\ : SLE
      port map(D => \waddr_gray[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[15]_net_1\);
    
    \wsync2_rptr[5]\ : SLE
      port map(D => \wsync1_rptr[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[5]_net_1\);
    
    \rgraynext[22]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIN3U66_S[23]\, B => 
        \rbinaddr_RNIPCKS5_S[22]\, Y => \rgraynext[22]_net_1\);
    
    \rbinaddr[5]\ : SLE
      port map(D => \rbinaddr_3[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[5]_net_1\);
    
    \raddr_gray[20]\ : SLE
      port map(D => \rgraynext[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[20]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_70\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIMR7H6_S[24]\, B => 
        \rsync2_wptr[23]_net_1\, C => \rbinaddr_RNIN3U66_S[23]\, 
        Y => fifo_empty_xhdl3_0_N_26);
    
    \wsync1_rptr[17]\ : SLE
      port map(D => \raddr_gray[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[17]_net_1\);
    
    \wbinaddr[10]\ : SLE
      port map(D => \wbinaddr_2[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[10]_net_1\);
    
    un13_writefull_0_I_69 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[23]_net_1\, B => 
        \wgraynext[22]_net_1\, C => \wgraynext[23]_net_1\, D => 
        \wsync2_rptr[22]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[10]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[11]\);
    
    \rgraynext[28]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI03P48_S[29]\, B => 
        \rbinaddr_RNIS5FQ7_S[28]\, Y => \rgraynext[28]_net_1\);
    
    \wgraynext[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI3T3D2_S[12]\, B => 
        \wbinaddr_RNI2I612_S[11]\, Y => \wgraynext[11]_net_1\);
    
    un13_writefull_0_I_63 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[21]_net_1\, B => 
        \wgraynext[20]_net_1\, C => \wgraynext[21]_net_1\, D => 
        \wsync2_rptr[20]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[9]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[10]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_75\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[2]_net_1\, B => 
        \rbinaddr_RNIB21T_S[2]\, C => \rbinaddr_RNINNN01_S[3]\, D
         => fifo_empty_xhdl3_0_N_21, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[0]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[1]\);
    
    \wgraynext[13]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI8MU43_S[14]\, B => 
        \wbinaddr_RNI591P2_S[13]\, Y => \wgraynext[13]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[9]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIKD0N1_S[9]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[9]\);
    
    \waddr_gray[28]\ : SLE
      port map(D => \wgraynext[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[28]_net_1\);
    
    \raddr_gray[32]\ : SLE
      port map(D => \rbinaddr_RNIN7P39_S[32]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[32]_net_1\);
    
    \wsync2_rptr[28]\ : SLE
      port map(D => \wsync1_rptr[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[28]_net_1\);
    
    \rbinaddr[20]\ : SLE
      port map(D => \rbinaddr_3[20]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[20]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_28\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI02185_S[20]\, B => 
        \rsync2_wptr[19]_net_1\, C => \rbinaddr_RNI5ENT4_S[19]\, 
        Y => fifo_empty_xhdl3_0_N_61);
    
    \wsync1_rptr[4]\ : SLE
      port map(D => \raddr_gray[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[4]_net_1\);
    
    un13_writefull_0_I_45 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[15]_net_1\, B => 
        \wgraynext[14]_net_1\, C => \wgraynext[15]\, D => 
        \wsync2_rptr[14]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[6]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[7]\);
    
    \rsync1_wptr[32]\ : SLE
      port map(D => \waddr_gray[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[32]_net_1\);
    
    \rbinaddr[4]\ : SLE
      port map(D => \rbinaddr_3[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[4]_net_1\);
    
    \rsync2_wptr[14]\ : SLE
      port map(D => \rsync1_wptr[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[14]_net_1\);
    
    \rsync2_wptr[6]\ : SLE
      port map(D => \rsync1_wptr[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[6]_net_1\);
    
    \rsync1_wptr[19]\ : SLE
      port map(D => \waddr_gray[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[19]_net_1\);
    
    \rbinaddr[23]\ : SLE
      port map(D => \rbinaddr_3[23]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[23]_net_1\);
    
    un13_writefull_0_I_81 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[27]_net_1\, B => 
        \wgraynext[26]_net_1\, C => \wgraynext[27]_net_1\, D => 
        \wsync2_rptr[26]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[12]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[13]\);
    
    \rsync2_wptr[10]\ : SLE
      port map(D => \rsync1_wptr[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[10]_net_1\);
    
    \rsync1_wptr[0]\ : SLE
      port map(D => \waddr_gray[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[0]_net_1\);
    
    \wsync2_rptr[25]\ : SLE
      port map(D => \wsync1_rptr[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[25]_net_1\);
    
    \wbinaddr[15]\ : SLE
      port map(D => \wbinaddr_2[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[15]_net_1\);
    
    \rgraynext[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIHNIF1_S[7]\, B => 
        \rbinaddr_RNI1URB1_S[6]\, Y => \rgraynext[6]_net_1\);
    
    un13_writefull_0_I_46_1 : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIHJPS3_S[16]\, B => 
        \wbinaddr_RNIC4SG3_S[15]\, Y => \wgraynext[15]\);
    
    \Read_Bin_Ptr.rbinaddr_3[17]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI0P594_S[17]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[17]\);
    
    \rsync1_wptr[5]\ : SLE
      port map(D => \waddr_gray[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[5]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[22]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI9BD46_S[22]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[22]\);
    
    \rsync2_wptr[21]\ : SLE
      port map(D => \rsync1_wptr[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[21]_net_1\);
    
    \wbinaddr_RNICPBG6[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_22, S
         => \wbinaddr_RNICPBG6_S[23]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_23);
    
    \waddr_gray[25]\ : SLE
      port map(D => \wgraynext[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[25]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[23]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNICPBG6_S[23]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[23]\);
    
    \rbinaddr[1]\ : SLE
      port map(D => \rbinaddr_3[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[1]_net_1\);
    
    \raddr_gray[14]\ : SLE
      port map(D => \rgraynext[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[14]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_27\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[18]_net_1\, B => 
        \rbinaddr_RNI2JEJ4_S[18]\, C => \rbinaddr_RNI5ENT4_S[19]\, 
        D => fifo_empty_xhdl3_0_N_61, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[8]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[9]\);
    
    \wsync2_rptr[22]\ : SLE
      port map(D => \wsync1_rptr[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[22]_net_1\);
    
    \wsync1_rptr[24]\ : SLE
      port map(D => \raddr_gray[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[24]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[1]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI7E1J_S[1]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[1]\);
    
    un13_writefull_0_I_9 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[3]_net_1\, B => 
        \wgraynext[2]_net_1\, C => \wgraynext[3]_net_1\, D => 
        \wsync2_rptr[2]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[0]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[1]\);
    
    \rsync1_wptr[13]\ : SLE
      port map(D => \waddr_gray[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[13]_net_1\);
    
    \rbinaddr[16]\ : SLE
      port map(D => \rbinaddr_3[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[16]_net_1\);
    
    \wbinaddr[32]\ : SLE
      port map(D => \wbinaddr_2[32]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[32]_net_1\);
    
    \waddr_gray[13]\ : SLE
      port map(D => \wgraynext[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[13]_net_1\);
    
    \rsync1_wptr[21]\ : SLE
      port map(D => \waddr_gray[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[21]_net_1\);
    
    \rbinaddr_RNIPFEP8[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[31]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_30, S
         => \rbinaddr_RNIPFEP8_S[31]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_31);
    
    \rsync1_wptr[14]\ : SLE
      port map(D => \waddr_gray[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[14]_net_1\);
    
    \wsync2_rptr[18]\ : SLE
      port map(D => \wsync1_rptr[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[18]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[24]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIG8AS6_S[24]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[24]\);
    
    \Write_Bin_Ptr.wbinaddr_2[19]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI67I05_S[19]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[19]\);
    
    \rbinaddr_RNIP95G7[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_26, S
         => \rbinaddr_RNIP95G7_S[27]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_27);
    
    \rbinaddr[7]\ : SLE
      port map(D => \rbinaddr_3[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[7]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[20]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI6IGC5_S[20]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[20]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_33\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[24]_net_1\, B => 
        \rbinaddr_RNIMR7H6_S[24]\, C => \rbinaddr_RNIMKHR6_S[25]\, 
        D => fifo_empty_xhdl3_0_N_56, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[11]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[12]\);
    
    \wbinaddr_RNIHJPS3[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_15, S
         => \wbinaddr_RNIHJPS3_S[16]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_16);
    
    \rgraynext[24]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIMKHR6_S[25]\, B => 
        \rbinaddr_RNIMR7H6_S[24]\, Y => \rgraynext[24]_net_1\);
    
    \raddr_gray[16]\ : SLE
      port map(D => \rgraynext[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[16]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \wbinaddr_RNI8MU43[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_13, S
         => \wbinaddr_RNI8MU43_S[14]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_14);
    
    \wgraynext[21]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI9BD46_S[22]\, B => 
        \wbinaddr_RNI7UEO5_S[21]\, Y => \wgraynext[21]_net_1\);
    
    \waddr_gray[24]\ : SLE
      port map(D => \wgraynext[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[24]_net_1\);
    
    \waddr_gray[1]\ : SLE
      port map(D => \wgraynext[1]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[1]_net_1\);
    
    \wsync2_rptr[15]\ : SLE
      port map(D => \wsync1_rptr[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[15]_net_1\);
    
    \wgraynext[23]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIG8AS6_S[24]\, B => 
        \wbinaddr_RNICPBG6_S[23]\, Y => \wgraynext[23]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[7]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIM4P31_S[7]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[7]\);
    
    \wbinaddr_RNI591P2[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_12, S
         => \wbinaddr_RNI591P2_S[13]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_13);
    
    \wbinaddr_RNI7UEO5[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_20, S
         => \wbinaddr_RNI7UEO5_S[21]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_21);
    
    \wsync2_rptr[12]\ : SLE
      port map(D => \wsync1_rptr[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[12]_net_1\);
    
    \wsync1_rptr[14]\ : SLE
      port map(D => \raddr_gray[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[14]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[2]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNINKQL_S[2]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[2]\);
    
    \wbinaddr_RNIPD1S9[32]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[32]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_31, S
         => \wbinaddr_RNIPD1S9_S[32]\, Y => OPEN, FCO => OPEN);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_39\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[12]_net_1\, B => 
        \rbinaddr_RNI56QL2_S[12]\, C => \rbinaddr_RNI2R203_S[13]\, 
        D => fifo_empty_xhdl3_0_N_51, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[5]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[6]\);
    
    \Read_Bin_Ptr.rbinaddr_3[8]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI2I9J1_S[8]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[8]\);
    
    \wsync1_rptr[5]\ : SLE
      port map(D => \raddr_gray[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[5]_net_1\);
    
    \wbinaddr_RNIMU1G9[31]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[31]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_30, S
         => \wbinaddr_RNIMU1G9_S[31]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_31);
    
    \rsync1_wptr[1]\ : SLE
      port map(D => \waddr_gray[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[1]_net_1\);
    
    \wgraynext[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI591P2_S[13]\, B => 
        \wbinaddr_RNI3T3D2_S[12]\, Y => \wgraynext[12]_net_1\);
    
    \wbinaddr[27]\ : SLE
      port map(D => \wbinaddr_2[27]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[27]_net_1\);
    
    \rgraynext[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNII5581_S[5]\, B => 
        \rbinaddr_RNI4EE41_S[4]\, Y => \rgraynext[4]_net_1\);
    
    \wsync2_rptr[2]\ : SLE
      port map(D => \wsync1_rptr[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[2]_net_1\);
    
    \wgraynext[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIMU1G9_S[31]\, B => 
        \wbinaddr_RNIKG249_S[30]\, Y => \wgraynext[30]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[26]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIR97K7_S[26]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[26]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_40\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI0HBA3_S[14]\, B => 
        \rsync2_wptr[13]_net_1\, C => \rbinaddr_RNI2R203_S[13]\, 
        Y => fifo_empty_xhdl3_0_N_51);
    
    \wbinaddr_RNIC4SG3[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_14, S
         => \wbinaddr_RNIC4SG3_S[15]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_15);
    
    \raddr_gray[1]\ : SLE
      port map(D => \rgraynext[1]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[1]_net_1\);
    
    \rsync1_wptr[27]\ : SLE
      port map(D => \waddr_gray[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[27]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_94\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI1URB1_S[6]\, B => 
        \rsync2_wptr[5]_net_1\, C => \rbinaddr_RNII5581_S[5]\, Y
         => fifo_empty_xhdl3_0_N_6);
    
    \rsync2_wptr[13]\ : SLE
      port map(D => \rsync1_wptr[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[13]_net_1\);
    
    \raddr_gray[31]\ : SLE
      port map(D => \rgraynext[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[31]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_45\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[14]_net_1\, B => 
        \rbinaddr_RNI0HBA3_S[14]\, C => \rbinaddr_RNIV7KK3_S[15]\, 
        D => fifo_empty_xhdl3_0_N_46, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[6]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[7]\);
    
    \wbinaddr[19]\ : SLE
      port map(D => \wbinaddr_2[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[19]_net_1\);
    
    \rsync1_wptr[20]\ : SLE
      port map(D => \waddr_gray[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[20]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_10\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIN7P39_S[32]\, B => 
        \rsync2_wptr[31]_net_1\, C => \rbinaddr_RNIPFEP8_S[31]\, 
        Y => fifo_empty_xhdl3_0_N_76);
    
    \rsync2_wptr[22]\ : SLE
      port map(D => \rsync1_wptr[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[22]_net_1\);
    
    un13_writefull_0_I_15 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[5]_net_1\, B => 
        \wgraynext[4]_net_1\, C => \wgraynext[5]_net_1\, D => 
        \wsync2_rptr[4]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[1]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[2]\);
    
    \wbinaddr_RNICHI61[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_7, S
         => \wbinaddr_RNICHI61_S[8]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_8);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_81\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[8]_net_1\, B => 
        \rbinaddr_RNI2I9J1_S[8]\, C => \rbinaddr_RNIKD0N1_S[9]\, 
        D => fifo_empty_xhdl3_0_N_16, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[3]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[4]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_15\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[28]_net_1\, B => 
        \rbinaddr_RNIS5FQ7_S[28]\, C => \rbinaddr_RNI03P48_S[29]\, 
        D => fifo_empty_xhdl3_0_N_71, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[13]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[14]\);
    
    \wsync1_rptr[20]\ : SLE
      port map(D => \raddr_gray[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[20]_net_1\);
    
    \wsync1_rptr[29]\ : SLE
      port map(D => \raddr_gray[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[29]_net_1\);
    
    un13_writefull_0_I_39 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[13]_net_1\, B => 
        \wgraynext[12]_net_1\, C => \wgraynext[13]_net_1\, D => 
        \wsync2_rptr[12]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[5]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[6]\);
    
    \rbinaddr[0]\ : SLE
      port map(D => \rbinaddr_3[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[0]_net_1\);
    
    un13_writefull_0_I_33 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[11]_net_1\, B => 
        \wgraynext[10]_net_1\, C => \wgraynext[11]_net_1\, D => 
        \wsync2_rptr[10]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[4]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[5]\);
    
    \rsync2_wptr[30]\ : SLE
      port map(D => \rsync1_wptr[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[30]_net_1\);
    
    \rsync1_wptr[26]\ : SLE
      port map(D => \waddr_gray[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[26]_net_1\);
    
    \wbinaddr_RNI2I612[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_10, S
         => \wbinaddr_RNI2I612_S[11]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_11);
    
    \raddr_gray[17]\ : SLE
      port map(D => \rgraynext[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[17]_net_1\);
    
    \rbinaddr[25]\ : SLE
      port map(D => \rbinaddr_3[25]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[25]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[17]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIN3N84_S[17]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[17]\);
    
    un9_writefull : CFG4
      generic map(INIT => x"0220")

      port map(A => \un7_writefull\, B => un13_writefull_0_N_2, C
         => \wsync2_rptr[32]_net_1\, D => 
        \wbinaddr_RNIPD1S9_S[32]\, Y => un9_writefull_0);
    
    \rsync2_wptr[17]\ : SLE
      port map(D => \rsync1_wptr[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[17]_net_1\);
    
    \rbinaddr_RNIB21T[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_1, S
         => \rbinaddr_RNIB21T_S[2]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_2);
    
    \Write_Bin_Ptr.wbinaddr_2[4]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIQ4DR_S[4]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[4]\);
    
    \wbinaddr_RNIO88G[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_0_cy, 
        S => \wbinaddr_RNIO88G_S[0]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_0);
    
    \wsync2_rptr[6]\ : SLE
      port map(D => \wsync1_rptr[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[6]_net_1\);
    
    \wsync1_rptr[28]\ : SLE
      port map(D => \raddr_gray[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[28]_net_1\);
    
    \rgraynext[16]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0P594_S[17]\, B => 
        \rbinaddr_RNIVVSU3_S[16]\, Y => \rgraynext[16]_net_1\);
    
    \rgraynext[19]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI02185_S[20]\, B => 
        \rbinaddr_RNI5ENT4_S[19]\, Y => \rgraynext[19]_net_1\);
    
    \wsync2_rptr[26]\ : SLE
      port map(D => \wsync1_rptr[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[26]_net_1\);
    
    \wgraynext[22]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNICPBG6_S[23]\, B => 
        \wbinaddr_RNI9BD46_S[22]\, Y => \wgraynext[22]_net_1\);
    
    \wgraynext[14]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIC4SG3_S[15]\, B => 
        \wbinaddr_RNI8MU43_S[14]\, Y => \wgraynext[14]_net_1\);
    
    \waddr_gray[4]\ : SLE
      port map(D => \wgraynext[4]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[4]_net_1\);
    
    \rgraynext[17]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI2JEJ4_S[18]\, B => 
        \rbinaddr_RNI0P594_S[17]\, Y => \rgraynext[17]_net_1\);
    
    \raddr_gray[24]\ : SLE
      port map(D => \rgraynext[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[24]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[6]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI1URB1_S[6]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[6]\);
    
    \rbinaddr_RNI2JEJ4[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_17, S
         => \rbinaddr_RNI2JEJ4_S[18]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_18);
    
    \waddr_gray[23]\ : SLE
      port map(D => \wgraynext[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[23]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[5]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIDE6U_S[5]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[5]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \rgraynext[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI1URB1_S[6]\, B => 
        \rbinaddr_RNII5581_S[5]\, Y => \rgraynext[5]_net_1\);
    
    \wsync1_rptr[10]\ : SLE
      port map(D => \raddr_gray[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[10]_net_1\);
    
    \wgraynext[28]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIJ33O8_S[29]\, B => 
        \wbinaddr_RNIAF4C8_S[28]\, Y => \wgraynext[28]_net_1\);
    
    \rbinaddr[28]\ : SLE
      port map(D => \rbinaddr_3[28]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[28]_net_1\);
    
    \wbinaddr[26]\ : SLE
      port map(D => \wbinaddr_2[26]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[26]_net_1\);
    
    \wsync1_rptr[19]\ : SLE
      port map(D => \raddr_gray[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[19]_net_1\);
    
    \wbinaddr[11]\ : SLE
      port map(D => \wbinaddr_2[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[11]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[32]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIN7P39_S[32]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[32]\);
    
    \rbinaddr_RNIMR7H6[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_23, S
         => \rbinaddr_RNIMR7H6_S[24]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_24);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_88\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI2I9J1_S[8]\, B => 
        \rsync2_wptr[7]_net_1\, C => \rbinaddr_RNIHNIF1_S[7]\, Y
         => fifo_empty_xhdl3_0_N_11);
    
    \wgraynext[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNICHI61_S[8]\, B => 
        \wbinaddr_RNIM4P31_S[7]\, Y => \wgraynext[7]_net_1\);
    
    un7_writefull : CFG2
      generic map(INIT => x"6")

      port map(A => \wgraynext[31]_net_1\, B => 
        \wsync2_rptr[31]_net_1\, Y => \un7_writefull\);
    
    \wgraynext[31]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIPD1S9_S[32]\, B => 
        \wbinaddr_RNIMU1G9_S[31]\, Y => \wgraynext[31]_net_1\);
    
    \wbinaddr_RNI6IGC5[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_19, S
         => \wbinaddr_RNI6IGC5_S[20]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_20);
    
    \wbinaddr[24]\ : SLE
      port map(D => \wbinaddr_2[24]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[24]_net_1\);
    
    \rbinaddr[21]\ : SLE
      port map(D => \rbinaddr_3[21]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[21]_net_1\);
    
    \raddr_gray[26]\ : SLE
      port map(D => \rgraynext[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[26]_net_1\);
    
    \wsync2_rptr[1]\ : SLE
      port map(D => \wsync1_rptr[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[1]_net_1\);
    
    \rsync1_wptr[22]\ : SLE
      port map(D => \waddr_gray[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[22]_net_1\);
    
    \rbinaddr[3]\ : SLE
      port map(D => \rbinaddr_3[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[3]_net_1\);
    
    \rsync2_wptr[9]\ : SLE
      port map(D => \rsync1_wptr[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[9]_net_1\);
    
    \rbinaddr[30]\ : SLE
      port map(D => \rbinaddr_3[30]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[30]_net_1\);
    
    \rsync2_wptr[7]\ : SLE
      port map(D => \rsync1_wptr[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[7]_net_1\);
    
    \rsync1_wptr[8]\ : SLE
      port map(D => \waddr_gray[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[8]_net_1\);
    
    \wsync1_rptr[18]\ : SLE
      port map(D => \raddr_gray[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[18]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[8]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNICHI61_S[8]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[8]\);
    
    \rbinaddr[9]\ : SLE
      port map(D => \rbinaddr_3[9]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[9]_net_1\);
    
    \waddr_gray[30]\ : SLE
      port map(D => \wgraynext[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[30]_net_1\);
    
    un13_writefull_0_I_58_1 : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI6IGC5_S[20]\, B => 
        \wbinaddr_RNI67I05_S[19]\, Y => \wgraynext[19]\);
    
    \wbinaddr[6]\ : SLE
      port map(D => \wbinaddr_2[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[6]_net_1\);
    
    \wsync2_rptr[16]\ : SLE
      port map(D => \wsync1_rptr[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[16]_net_1\);
    
    \waddr_gray[11]\ : SLE
      port map(D => \wgraynext[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[11]_net_1\);
    
    \rsync2_wptr[16]\ : SLE
      port map(D => \rsync1_wptr[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[16]_net_1\);
    
    \wsync2_rptr[32]\ : SLE
      port map(D => \wsync1_rptr[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[32]_net_1\);
    
    \wsync1_rptr[2]\ : SLE
      port map(D => \raddr_gray[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[2]_net_1\);
    
    \raddr_gray[4]\ : SLE
      port map(D => \rgraynext[4]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[4]_net_1\);
    
    \rsync2_wptr[2]\ : SLE
      port map(D => \rsync1_wptr[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[2]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[28]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIS5FQ7_S[28]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[28]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_87\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[6]_net_1\, B => 
        \rbinaddr_RNI1URB1_S[6]\, C => \rbinaddr_RNIHNIF1_S[7]\, 
        D => fifo_empty_xhdl3_0_N_11, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[2]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[3]\);
    
    \rbinaddr[12]\ : SLE
      port map(D => \rbinaddr_3[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[12]_net_1\);
    
    \wsync2_rptr[21]\ : SLE
      port map(D => \wsync1_rptr[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[21]_net_1\);
    
    \wgraynext[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNINKQL_S[2]\, B => 
        \wbinaddr_RNI8SJO_S[3]\, Y => \wgraynext[2]_net_1\);
    
    \rsync2_wptr[29]\ : SLE
      port map(D => \rsync1_wptr[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[29]_net_1\);
    
    \wsync2_rptr[9]\ : SLE
      port map(D => \wsync1_rptr[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[9]_net_1\);
    
    \wgraynext[24]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNILO887_S[25]\, B => 
        \wbinaddr_RNIG8AS6_S[24]\, Y => \wgraynext[24]_net_1\);
    
    \rbinaddr[24]\ : SLE
      port map(D => \rbinaddr_3[24]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[24]_net_1\);
    
    \waddr_gray[5]\ : SLE
      port map(D => \wgraynext[5]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[5]_net_1\);
    
    un13_writefull_0_I_87 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[29]_net_1\, B => 
        \wgraynext[28]_net_1\, C => \wgraynext[29]_net_1\, D => 
        \wsync2_rptr[28]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[13]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[14]\);
    
    \wbinaddr_RNIN3N84[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_16, S
         => \wbinaddr_RNIN3N84_S[17]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_17);
    
    \wsync2_rptr[20]\ : SLE
      port map(D => \wsync1_rptr[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[20]_net_1\);
    
    \rsync2_wptr[25]\ : SLE
      port map(D => \rsync1_wptr[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[25]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_4\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIB21T_S[2]\, B => 
        \rsync2_wptr[1]_net_1\, C => \rbinaddr_RNI0EAP_S[1]\, Y
         => fifo_empty_xhdl3_0_N_81);
    
    \wbinaddr[23]\ : SLE
      port map(D => \wbinaddr_2[23]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[23]_net_1\);
    
    \waddr_gray[32]\ : SLE
      port map(D => \wbinaddr_RNIPD1S9_S[32]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[32]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_63\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[20]_net_1\, B => 
        \rbinaddr_RNI02185_S[20]\, C => \rbinaddr_RNISMAI5_S[21]\, 
        D => fifo_empty_xhdl3_0_N_31, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[9]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[10]\);
    
    \wbinaddr_RNIG8AS6[24]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[24]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_23, S
         => \wbinaddr_RNIG8AS6_S[24]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_24);
    
    \rsync1_wptr[6]\ : SLE
      port map(D => \waddr_gray[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[6]_net_1\);
    
    \rsync1_wptr[18]\ : SLE
      port map(D => \waddr_gray[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[18]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_22\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIS5FQ7_S[28]\, B => 
        \rsync2_wptr[27]_net_1\, C => \rbinaddr_RNIP95G7_S[27]\, 
        Y => fifo_empty_xhdl3_0_N_66);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_1\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[0]_net_1\, B => 
        \rbinaddr_RNIMQJL_S[0]\, C => \rbinaddr_RNI0EAP_S[1]\, D
         => fifo_empty_xhdl3_0_N_81, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \fifo_empty_xhdl3_0_data_tmp[0]\);
    
    \Write_Bin_Ptr.wbinaddr_2[11]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI2I612_S[11]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[11]\);
    
    \rgraynext[26]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIP95G7_S[27]\, B => 
        \rbinaddr_RNINER57_S[26]\, Y => \rgraynext[26]_net_1\);
    
    \rgraynext[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNISO3F8_S[30]\, B => 
        \rbinaddr_RNI03P48_S[29]\, Y => \rgraynext[29]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[9]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI3VB91_S[9]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[9]\);
    
    fifo_empty_xhdl3_RNO : CFG1
      generic map(INIT => "01")

      port map(A => fifo_empty_xhdl3_0_N_2, Y => 
        fifo_empty_xhdl3_0_N_2_i);
    
    \wsync1_rptr[6]\ : SLE
      port map(D => \raddr_gray[6]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[6]_net_1\);
    
    \rgraynext[27]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIS5FQ7_S[28]\, B => 
        \rbinaddr_RNIP95G7_S[27]\, Y => \rgraynext[27]_net_1\);
    
    \wsync2_rptr[11]\ : SLE
      port map(D => \wsync1_rptr[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[11]_net_1\);
    
    \raddr_gray[27]\ : SLE
      port map(D => \rgraynext[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[27]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[29]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIJ33O8_S[29]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[29]\);
    
    \rsync2_wptr[3]\ : SLE
      port map(D => \rsync1_wptr[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[3]_net_1\);
    
    \wsync2_rptr[23]\ : SLE
      port map(D => \wsync1_rptr[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[23]_net_1\);
    
    \wbinaddr_RNIR97K7[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_25, S
         => \wbinaddr_RNIR97K7_S[26]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_26);
    
    \rsync1_wptr[25]\ : SLE
      port map(D => \waddr_gray[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[25]_net_1\);
    
    \raddr_gray[5]\ : SLE
      port map(D => \rgraynext[5]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[5]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_69\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[22]_net_1\, B => 
        \rbinaddr_RNIPCKS5_S[22]\, C => \rbinaddr_RNIN3U66_S[23]\, 
        D => fifo_empty_xhdl3_0_N_26, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[10]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[11]\);
    
    un13_writefull_0_I_75 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[25]_net_1\, B => 
        \wgraynext[24]_net_1\, C => \wgraynext[25]_net_1\, D => 
        \wsync2_rptr[24]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[11]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[12]\);
    
    \Read_Bin_Ptr.rbinaddr_3[22]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIPCKS5_S[22]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[22]\);
    
    \wbinaddr[12]\ : SLE
      port map(D => \wbinaddr_2[12]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[12]_net_1\);
    
    \rbinaddr_RNINNN01[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_2, S
         => \rbinaddr_RNINNN01_S[3]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_3);
    
    \raddr_gray[19]\ : SLE
      port map(D => \rgraynext[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[19]_net_1\);
    
    \wsync2_rptr[10]\ : SLE
      port map(D => \wsync1_rptr[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[10]_net_1\);
    
    \wsync2_rptr[24]\ : SLE
      port map(D => \wsync1_rptr[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[24]_net_1\);
    
    \wbinaddr[20]\ : SLE
      port map(D => \wbinaddr_2[20]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[20]_net_1\);
    
    \wbinaddr_RNILO887[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_24, S
         => \wbinaddr_RNILO887_S[25]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_25);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_34\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNINER57_S[26]\, B => 
        \rsync2_wptr[25]_net_1\, C => \rbinaddr_RNIMKHR6_S[25]\, 
        Y => fifo_empty_xhdl3_0_N_56);
    
    \raddr_gray[30]\ : SLE
      port map(D => \rgraynext[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[30]_net_1\);
    
    \wgraynext[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI1PV01_S[6]\, B => 
        \wbinaddr_RNIDE6U_S[5]\, Y => \wgraynext[5]_net_1\);
    
    \raddr_gray[12]\ : SLE
      port map(D => \rgraynext[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[12]_net_1\);
    
    \wsync1_rptr[30]\ : SLE
      port map(D => \raddr_gray[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[30]_net_1\);
    
    \wsync1_rptr[1]\ : SLE
      port map(D => \raddr_gray[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[1]_net_1\);
    
    \rbinaddr_RNI1URB1[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_5, S
         => \rbinaddr_RNI1URB1_S[6]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_6);
    
    fifo_empty_xhdl3 : SLE
      port map(D => fifo_empty_xhdl3_0_N_2_i, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rdch_fifo_empty\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_9\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[30]_net_1\, B => 
        \rbinaddr_RNISO3F8_S[30]\, C => \rbinaddr_RNIPFEP8_S[31]\, 
        D => fifo_empty_xhdl3_0_N_76, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[14]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[15]\);
    
    \rsync2_wptr[4]\ : SLE
      port map(D => \rsync1_wptr[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[4]_net_1\);
    
    \rbinaddr_RNI2I9J1[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_7, S
         => \rbinaddr_RNI2I9J1_S[8]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_8);
    
    fifo_empty_xhdl3_RNID8TH : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => \rdch_fifo_empty\, C => 
        rdch_fifo_rd_en_r, D => GND_net_1, FCI => VCC_net_1, S
         => OPEN, Y => OPEN, FCO => un3_rbinnext_cry_0_cy);
    
    \rsync2_wptr[24]\ : SLE
      port map(D => \rsync1_wptr[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[24]_net_1\);
    
    \wsync2_rptr[13]\ : SLE
      port map(D => \wsync1_rptr[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[13]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[31]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIMU1G9_S[31]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[31]\);
    
    un13_writefull_0_I_51 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[17]_net_1\, B => \wgraynext[16]\, 
        C => \wgraynext[17]\, D => \wsync2_rptr[16]_net_1\, FCI
         => \un13_writefull_0_data_tmp[7]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[8]\);
    
    \rsync1_wptr[29]\ : SLE
      port map(D => \waddr_gray[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[29]_net_1\);
    
    \rsync2_wptr[20]\ : SLE
      port map(D => \rsync1_wptr[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[20]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[2]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIB21T_S[2]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[2]\);
    
    \wbinaddr[25]\ : SLE
      port map(D => \wbinaddr_2[25]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[25]_net_1\);
    
    \rgraynext[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI4EE41_S[4]\, B => 
        \rbinaddr_RNINNN01_S[3]\, Y => \rgraynext[3]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[4]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI4EE41_S[4]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[4]\);
    
    \wsync2_rptr[14]\ : SLE
      port map(D => \wsync1_rptr[14]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[14]_net_1\);
    
    un13_writefull_0_I_53_1 : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIN3N84_S[17]\, B => 
        \wbinaddr_RNIHJPS3_S[16]\, Y => \wgraynext[16]\);
    
    \rgraynext[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0EAP_S[1]\, B => 
        \rbinaddr_RNIMQJL_S[0]\, Y => \rgraynext[0]_net_1\);
    
    \waddr_gray[7]\ : SLE
      port map(D => \wgraynext[7]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[7]_net_1\);
    
    \waddr_gray[21]\ : SLE
      port map(D => \wgraynext[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[21]_net_1\);
    
    \rgraynext[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIB21T_S[2]\, B => 
        \rbinaddr_RNI0EAP_S[1]\, Y => \rgraynext[1]_net_1\);
    
    un13_writefull_0_I_21 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[7]_net_1\, B => 
        \wgraynext[6]_net_1\, C => \wgraynext[7]_net_1\, D => 
        \wsync2_rptr[6]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[2]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[3]\);
    
    \rgraynext[30]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIPFEP8_S[31]\, B => 
        \rbinaddr_RNISO3F8_S[30]\, Y => \rgraynext[30]_net_1\);
    
    \waddr_gray[9]\ : SLE
      port map(D => \wgraynext[9]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[9]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[18]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI2JEJ4_S[18]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[18]\);
    
    \wbinaddr_RNI289L1[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_9, S
         => \wbinaddr_RNI289L1_S[10]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_10);
    
    \rsync1_wptr[23]\ : SLE
      port map(D => \waddr_gray[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[23]_net_1\);
    
    \wsync1_rptr[9]\ : SLE
      port map(D => \raddr_gray[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[9]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[24]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIMR7H6_S[24]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[24]\);
    
    \rbinaddr[26]\ : SLE
      port map(D => \rbinaddr_3[26]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[26]_net_1\);
    
    \wbinaddr[8]\ : SLE
      port map(D => \wbinaddr_2[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[8]_net_1\);
    
    \rsync1_wptr[24]\ : SLE
      port map(D => \waddr_gray[24]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[24]_net_1\);
    
    \rgraynext[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIEV812_S[10]\, B => 
        \rbinaddr_RNIKD0N1_S[9]\, Y => \rgraynext[9]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[15]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIC4SG3_S[15]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[15]\);
    
    \Read_Bin_Ptr.rbinaddr_3[26]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNINER57_S[26]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[26]\);
    
    \rbinaddr_RNIN7P39[32]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[32]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_31, S
         => \rbinaddr_RNIN7P39_S[32]\, Y => OPEN, FCO => OPEN);
    
    \rbinaddr[19]\ : SLE
      port map(D => \rbinaddr_3[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[19]_net_1\);
    
    \waddr_gray[19]\ : SLE
      port map(D => \wgraynext[19]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[19]_net_1\);
    
    un13_writefull_0_I_59_1 : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI67I05_S[19]\, B => 
        \wbinaddr_RNIUKKK4_S[18]\, Y => \wgraynext[18]\);
    
    \wbinaddr[2]\ : SLE
      port map(D => \wbinaddr_2[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[2]_net_1\);
    
    \wsync2_rptr[0]\ : SLE
      port map(D => \wsync1_rptr[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[0]_net_1\);
    
    \rbinaddr[17]\ : SLE
      port map(D => \rbinaddr_3[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[17]_net_1\);
    
    \raddr_gray[18]\ : SLE
      port map(D => \rgraynext[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[18]_net_1\);
    
    \rbinaddr[31]\ : SLE
      port map(D => \rbinaddr_3[31]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[31]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[27]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI2S508_S[27]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[27]\);
    
    un13_writefull_0_I_52_1 : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIUKKK4_S[18]\, B => 
        \wbinaddr_RNIN3N84_S[17]\, Y => \wgraynext[17]\);
    
    \raddr_gray[7]\ : SLE
      port map(D => \rgraynext[7]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[7]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[0]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIO88G_S[0]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[0]\);
    
    \raddr_gray[9]\ : SLE
      port map(D => \rgraynext[9]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[9]_net_1\);
    
    \wbinaddr_RNI9BD46[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_21, S
         => \wbinaddr_RNI9BD46_S[22]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_22);
    
    \Read_Bin_Ptr.rbinaddr_3[31]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIPFEP8_S[31]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[31]\);
    
    \rbinaddr_RNI9IHB2[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_10, S
         => \rbinaddr_RNI9IHB2_S[11]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_11);
    
    \raddr_gray[13]\ : SLE
      port map(D => \rgraynext[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[13]_net_1\);
    
    \rbinaddr_RNI2R203[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_12, S
         => \rbinaddr_RNI2R203_S[13]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_13);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_51\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[10]_net_1\, B => 
        \rbinaddr_RNIEV812_S[10]\, C => \rbinaddr_RNI9IHB2_S[11]\, 
        D => fifo_empty_xhdl3_0_N_41, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[5]\);
    
    \wsync2_rptr[31]\ : SLE
      port map(D => \wsync1_rptr[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[31]_net_1\);
    
    \wbinaddr[18]\ : SLE
      port map(D => \wbinaddr_2[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[18]_net_1\);
    
    \rsync2_wptr[18]\ : SLE
      port map(D => \rsync1_wptr[18]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[18]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[30]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNISO3F8_S[30]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[30]\);
    
    \rbinaddr_RNIV7KK3[15]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[15]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_14, S
         => \rbinaddr_RNIV7KK3_S[15]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_15);
    
    \Read_Bin_Ptr.rbinaddr_3[23]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIN3U66_S[23]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[23]\);
    
    \rgraynext[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNINNN01_S[3]\, B => 
        \rbinaddr_RNIB21T_S[2]\, Y => \rgraynext[2]_net_1\);
    
    \raddr_gray[11]\ : SLE
      port map(D => \rgraynext[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[11]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[12]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI56QL2_S[12]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[12]\);
    
    \rbinaddr_RNIS5FQ7[28]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[28]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_27, S
         => \rbinaddr_RNIS5FQ7_S[28]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_28);
    
    \wsync2_rptr[30]\ : SLE
      port map(D => \wsync1_rptr[30]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[30]_net_1\);
    
    \raddr_gray[29]\ : SLE
      port map(D => \rgraynext[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[29]_net_1\);
    
    \rsync2_wptr[23]\ : SLE
      port map(D => \rsync1_wptr[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[23]_net_1\);
    
    \rgraynext[15]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIVVSU3_S[16]\, B => 
        \rbinaddr_RNIV7KK3_S[15]\, Y => \rgraynext[15]_net_1\);
    
    \wsync1_rptr[26]\ : SLE
      port map(D => \raddr_gray[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[26]_net_1\);
    
    \wbinaddr_RNIUKKK4[18]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[18]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_17, S
         => \wbinaddr_RNIUKKK4_S[18]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_18);
    
    \wbinaddr_RNI3VB91[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_8, S
         => \wbinaddr_RNI3VB91_S[9]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_9);
    
    \wbinaddr[29]\ : SLE
      port map(D => \wbinaddr_2[29]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[29]_net_1\);
    
    \rgraynext[31]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIN7P39_S[32]\, B => 
        \rbinaddr_RNIPFEP8_S[31]\, Y => \rgraynext[31]_net_1\);
    
    \raddr_gray[22]\ : SLE
      port map(D => \rgraynext[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[22]_net_1\);
    
    \wsync1_rptr[21]\ : SLE
      port map(D => \raddr_gray[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[21]_net_1\);
    
    \waddr_gray[17]\ : SLE
      port map(D => \wgraynext[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[17]_net_1\);
    
    \rsync1_wptr[9]\ : SLE
      port map(D => \waddr_gray[9]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[9]_net_1\);
    
    \rgraynext[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI9IHB2_S[11]\, B => 
        \rbinaddr_RNIEV812_S[10]\, Y => \rgraynext[10]_net_1\);
    
    \rbinaddr_RNISMAI5[21]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[21]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_20, S
         => \rbinaddr_RNISMAI5_S[21]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_21);
    
    fifo_full_xhdl2_RNIA4FD : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => \fifo_full_xhdl2\, C => 
        rdch_fifo_wr_en_r, D => GND_net_1, FCI => VCC_net_1, S
         => OPEN, Y => OPEN, FCO => un3_wbinnext_cry_0_cy);
    
    \wsync2_rptr[3]\ : SLE
      port map(D => \wsync1_rptr[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[3]_net_1\);
    
    \wbinaddr_RNIKG249[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_29, S
         => \wbinaddr_RNIKG249_S[30]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_30);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_82\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIEV812_S[10]\, B => 
        \rsync2_wptr[9]_net_1\, C => \rbinaddr_RNIKD0N1_S[9]\, Y
         => fifo_empty_xhdl3_0_N_16);
    
    \rsync1_wptr[7]\ : SLE
      port map(D => \waddr_gray[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[7]_net_1\);
    
    \rbinaddr_RNISO3F8[30]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[30]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_29, S
         => \rbinaddr_RNISO3F8_S[30]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_30);
    
    \rbinaddr[6]\ : SLE
      port map(D => \rbinaddr_3[6]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[6]_net_1\);
    
    \rbinaddr[10]\ : SLE
      port map(D => \rbinaddr_3[10]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[10]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[3]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI8SJO_S[3]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[3]\);
    
    \wgraynext[26]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI2S508_S[27]\, B => 
        \wbinaddr_RNIR97K7_S[26]\, Y => \wgraynext[26]_net_1\);
    
    \wgraynext[29]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIKG249_S[30]\, B => 
        \wbinaddr_RNIJ33O8_S[29]\, Y => \wgraynext[29]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_58\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI2JEJ4_S[18]\, B => 
        \rsync2_wptr[17]_net_1\, C => \rbinaddr_RNI0P594_S[17]\, 
        Y => fifo_empty_xhdl3_0_N_36);
    
    \wgraynext[27]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIAF4C8_S[28]\, B => 
        \wbinaddr_RNI2S508_S[27]\, Y => \wgraynext[27]_net_1\);
    
    \wsync2_rptr[29]\ : SLE
      port map(D => \wsync1_rptr[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[29]_net_1\);
    
    \rsync2_wptr[27]\ : SLE
      port map(D => \rsync1_wptr[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[27]_net_1\);
    
    \rsync1_wptr[2]\ : SLE
      port map(D => \waddr_gray[2]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[2]_net_1\);
    
    \rbinaddr[13]\ : SLE
      port map(D => \rbinaddr_3[13]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[13]_net_1\);
    
    \waddr_gray[6]\ : SLE
      port map(D => \wgraynext[6]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[6]_net_1\);
    
    \rsync2_wptr[11]\ : SLE
      port map(D => \rsync1_wptr[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[11]_net_1\);
    
    \wsync1_rptr[16]\ : SLE
      port map(D => \raddr_gray[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[16]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[25]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIMKHR6_S[25]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[25]\);
    
    \wsync1_rptr[11]\ : SLE
      port map(D => \raddr_gray[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[11]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[18]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIUKKK4_S[18]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[18]\);
    
    \wgraynext[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI7E1J_S[1]\, B => 
        \wbinaddr_RNIO88G_S[0]\, Y => \wgraynext[0]_net_1\);
    
    \wsync2_rptr[7]\ : SLE
      port map(D => \wsync1_rptr[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[7]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[14]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI0HBA3_S[14]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[14]\);
    
    \wsync1_rptr[22]\ : SLE
      port map(D => \raddr_gray[22]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[22]_net_1\);
    
    \rsync1_wptr[11]\ : SLE
      port map(D => \waddr_gray[11]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[11]_net_1\);
    
    \rbinaddr_RNIVVSU3[16]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[16]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_15, S
         => \rbinaddr_RNIVVSU3_S[16]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_16);
    
    \wsync1_rptr[0]\ : SLE
      port map(D => \raddr_gray[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[0]_net_1\);
    
    \wbinaddr_RNINKQL[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_1, S
         => \wbinaddr_RNINKQL_S[2]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_2);
    
    \wbinaddr[30]\ : SLE
      port map(D => \wbinaddr_2[30]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[30]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_57\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[16]_net_1\, B => 
        \rbinaddr_RNIVVSU3_S[16]\, C => \rbinaddr_RNI0P594_S[17]\, 
        D => fifo_empty_xhdl3_0_N_36, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[7]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[8]\);
    
    \Read_Bin_Ptr.rbinaddr_3[16]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIVVSU3_S[16]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[16]\);
    
    \rbinaddr_RNII5581[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_4, S
         => \rbinaddr_RNII5581_S[5]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_5);
    
    \wbinaddr_RNI2S508[27]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[27]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_26, S
         => \wbinaddr_RNI2S508_S[27]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_27);
    
    \wbinaddr[21]\ : SLE
      port map(D => \wbinaddr_2[21]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[21]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[21]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI7UEO5_S[21]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[21]\);
    
    \wbinaddr[5]\ : SLE
      port map(D => \wbinaddr_2[5]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[5]_net_1\);
    
    \waddr_gray[29]\ : SLE
      port map(D => \wgraynext[29]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[29]_net_1\);
    
    \rbinaddr_RNINER57[26]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[26]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_25, S
         => \rbinaddr_RNINER57_S[26]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_26);
    
    \wbinaddr_RNI7E1J[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_0, S
         => \wbinaddr_RNI7E1J_S[1]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_1);
    
    \rbinaddr_RNI4EE41[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_3, S
         => \rbinaddr_RNI4EE41_S[4]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_4);
    
    \wsync2_rptr[8]\ : SLE
      port map(D => \wsync1_rptr[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[8]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[29]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI03P48_S[29]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[29]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_64\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIPCKS5_S[22]\, B => 
        \rsync2_wptr[21]_net_1\, C => \rbinaddr_RNISMAI5_S[21]\, 
        Y => fifo_empty_xhdl3_0_N_31);
    
    \wsync2_rptr[19]\ : SLE
      port map(D => \wsync1_rptr[19]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[19]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[21]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNISMAI5_S[21]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[21]\);
    
    \wsync1_rptr[25]\ : SLE
      port map(D => \raddr_gray[25]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[25]_net_1\);
    
    \waddr_gray[8]\ : SLE
      port map(D => \wgraynext[8]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[8]_net_1\);
    
    \raddr_gray[28]\ : SLE
      port map(D => \rgraynext[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[28]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_76\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNI4EE41_S[4]\, B => 
        \rsync2_wptr[3]_net_1\, C => \rbinaddr_RNINNN01_S[3]\, Y
         => fifo_empty_xhdl3_0_N_21);
    
    \waddr_gray[10]\ : SLE
      port map(D => \wgraynext[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[10]_net_1\);
    
    \rgraynext[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI2I9J1_S[8]\, B => 
        \rbinaddr_RNIHNIF1_S[7]\, Y => \rgraynext[7]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[20]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI02185_S[20]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[20]\);
    
    \wsync1_rptr[23]\ : SLE
      port map(D => \raddr_gray[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[23]_net_1\);
    
    \wbinaddr_RNI1PV01[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_5, S
         => \wbinaddr_RNI1PV01_S[6]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_6);
    
    \raddr_gray[6]\ : SLE
      port map(D => \rgraynext[6]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[6]_net_1\);
    
    \wsync2_rptr[27]\ : SLE
      port map(D => \wsync1_rptr[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[27]_net_1\);
    
    \rsync2_wptr[26]\ : SLE
      port map(D => \rsync1_wptr[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[26]_net_1\);
    
    un13_writefull_0_I_1 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[1]_net_1\, B => 
        \wgraynext[0]_net_1\, C => \wgraynext[1]_net_1\, D => 
        \wsync2_rptr[0]_net_1\, FCI => GND_net_1, S => OPEN, Y
         => OPEN, FCO => \un13_writefull_0_data_tmp[0]\);
    
    \rsync1_wptr[3]\ : SLE
      port map(D => \waddr_gray[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[3]_net_1\);
    
    \waddr_gray[16]\ : SLE
      port map(D => \wgraynext[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[16]_net_1\);
    
    \wbinaddr[4]\ : SLE
      port map(D => \wbinaddr_2[4]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[4]_net_1\);
    
    \rgraynext[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI56QL2_S[12]\, B => 
        \rbinaddr_RNI9IHB2_S[11]\, Y => \rgraynext[11]_net_1\);
    
    \wsync1_rptr[12]\ : SLE
      port map(D => \raddr_gray[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[12]_net_1\);
    
    \rsync2_wptr[0]\ : SLE
      port map(D => \rsync1_wptr[0]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[0]_net_1\);
    
    \rgraynext[25]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNINER57_S[26]\, B => 
        \rbinaddr_RNIMKHR6_S[25]\, Y => \rgraynext[25]_net_1\);
    
    \raddr_gray[23]\ : SLE
      port map(D => \rgraynext[23]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[23]_net_1\);
    
    \rgraynext[13]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI0HBA3_S[14]\, B => 
        \rbinaddr_RNI2R203_S[13]\, Y => \rgraynext[13]_net_1\);
    
    \rbinaddr[22]\ : SLE
      port map(D => \rbinaddr_3[22]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[22]_net_1\);
    
    \wbinaddr_RNI8SJO[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_2, S
         => \wbinaddr_RNI8SJO_S[3]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_3);
    
    \rsync2_wptr[5]\ : SLE
      port map(D => \rsync1_wptr[5]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[5]_net_1\);
    
    \rbinaddr_RNIN3U66[23]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[23]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_22, S
         => \rbinaddr_RNIN3U66_S[23]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_23);
    
    \wbinaddr[17]\ : SLE
      port map(D => \wbinaddr_2[17]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[17]_net_1\);
    
    \rgraynext[20]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNISMAI5_S[21]\, B => 
        \rbinaddr_RNI02185_S[20]\, Y => \rgraynext[20]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[7]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIHNIF1_S[7]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[7]\);
    
    \rbinaddr_RNI02185[20]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[20]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_19, S
         => \rbinaddr_RNI02185_S[20]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_20);
    
    \wgraynext[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIQ4DR_S[4]\, B => 
        \wbinaddr_RNI8SJO_S[3]\, Y => \wgraynext[3]_net_1\);
    
    fifo_full_xhdl2 : SLE
      port map(D => un9_writefull_0, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_full_xhdl2\);
    
    \Read_Bin_Ptr.rbinaddr_3[13]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI2R203_S[13]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[13]\);
    
    \Write_Bin_Ptr.wbinaddr_2[12]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI3T3D2_S[12]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[12]\);
    
    un13_writefull_0_I_57 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[19]_net_1\, B => \wgraynext[18]\, 
        C => \wgraynext[19]\, D => \wsync2_rptr[18]_net_1\, FCI
         => \un13_writefull_0_data_tmp[8]\, S => OPEN, Y => OPEN, 
        FCO => \un13_writefull_0_data_tmp[9]\);
    
    \Read_Bin_Ptr.rbinaddr_3[3]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNINNN01_S[3]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[3]\);
    
    \raddr_gray[21]\ : SLE
      port map(D => \rgraynext[21]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[21]_net_1\);
    
    \raddr_gray[15]\ : SLE
      port map(D => \rgraynext[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[15]_net_1\);
    
    \wsync1_rptr[15]\ : SLE
      port map(D => \raddr_gray[15]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[15]_net_1\);
    
    \raddr_gray[8]\ : SLE
      port map(D => \rgraynext[8]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[8]_net_1\);
    
    \wsync1_rptr[3]\ : SLE
      port map(D => \raddr_gray[3]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[3]_net_1\);
    
    \wbinaddr[1]\ : SLE
      port map(D => \wbinaddr_2[1]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[1]_net_1\);
    
    \rsync1_wptr[17]\ : SLE
      port map(D => \waddr_gray[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[17]_net_1\);
    
    \waddr_gray[12]\ : SLE
      port map(D => \wgraynext[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[12]_net_1\);
    
    \wsync1_rptr[13]\ : SLE
      port map(D => \raddr_gray[13]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[13]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[13]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI591P2_S[13]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[13]\);
    
    \wsync2_rptr[17]\ : SLE
      port map(D => \wsync1_rptr[17]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[17]_net_1\);
    
    \rsync1_wptr[10]\ : SLE
      port map(D => \waddr_gray[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[10]_net_1\);
    
    \rsync2_wptr[12]\ : SLE
      port map(D => \rsync1_wptr[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[12]_net_1\);
    
    \rsync1_wptr[4]\ : SLE
      port map(D => \waddr_gray[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[4]_net_1\);
    
    \rbinaddr_RNIMKHR6[25]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[25]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_24, S
         => \rbinaddr_RNIMKHR6_S[25]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_25);
    
    \rbinaddr_RNI0HBA3[14]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[14]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_13, S
         => \rbinaddr_RNI0HBA3_S[14]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_14);
    
    \wbinaddr[7]\ : SLE
      port map(D => \wbinaddr_2[7]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[7]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[14]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI8MU43_S[14]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[14]\);
    
    un13_writefull_0_I_27 : ARI1
      generic map(INIT => x"68421")

      port map(A => \wsync2_rptr[9]_net_1\, B => 
        \wgraynext[8]_net_1\, C => \wgraynext[9]_net_1\, D => 
        \wsync2_rptr[8]_net_1\, FCI => 
        \un13_writefull_0_data_tmp[3]\, S => OPEN, Y => OPEN, FCO
         => \un13_writefull_0_data_tmp[4]\);
    
    \waddr_gray[27]\ : SLE
      port map(D => \wgraynext[27]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[27]_net_1\);
    
    \rsync1_wptr[28]\ : SLE
      port map(D => \waddr_gray[28]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[28]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[10]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI289L1_S[10]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[10]\);
    
    \wbinaddr_RNIM4P31[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_6, S
         => \wbinaddr_RNIM4P31_S[7]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_7);
    
    \wgraynext[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIDE6U_S[5]\, B => 
        \wbinaddr_RNIQ4DR_S[4]\, Y => \wgraynext[4]_net_1\);
    
    \wgraynext[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI7E1J_S[1]\, B => 
        \wbinaddr_RNINKQL_S[2]\, Y => \wgraynext[1]_net_1\);
    
    \rsync1_wptr[16]\ : SLE
      port map(D => \waddr_gray[16]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[16]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[5]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNII5581_S[5]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[5]\);
    
    \Write_Bin_Ptr.wbinaddr_2[25]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNILO887_S[25]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[25]\);
    
    \wbinaddr_RNIQ4DR[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_3, S
         => \wbinaddr_RNIQ4DR_S[4]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_4);
    
    \rbinaddr[8]\ : SLE
      port map(D => \rbinaddr_3[8]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[8]_net_1\);
    
    \rbinaddr[15]\ : SLE
      port map(D => \rbinaddr_3[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[15]_net_1\);
    
    \waddr_gray[2]\ : SLE
      port map(D => \wgraynext[2]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[2]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[0]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIMQJL_S[0]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[0]\);
    
    \rsync2_wptr[31]\ : SLE
      port map(D => \rsync1_wptr[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[31]_net_1\);
    
    \wsync1_rptr[7]\ : SLE
      port map(D => \raddr_gray[7]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[7]_net_1\);
    
    \rbinaddr_RNIPCKS5[22]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[22]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_21, S
         => \rbinaddr_RNIPCKS5_S[22]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_22);
    
    \wbinaddr[22]\ : SLE
      port map(D => \wbinaddr_2[22]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[22]_net_1\);
    
    \rsync2_wptr[1]\ : SLE
      port map(D => \rsync1_wptr[1]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync2_wptr[1]_net_1\);
    
    \raddr_gray[10]\ : SLE
      port map(D => \rgraynext[10]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[10]_net_1\);
    
    \rsync1_wptr[31]\ : SLE
      port map(D => \waddr_gray[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[31]_net_1\);
    
    \rgraynext[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIKD0N1_S[9]\, B => 
        \rbinaddr_RNI2I9J1_S[8]\, Y => \rgraynext[8]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[15]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIV7KK3_S[15]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[15]\);
    
    \rbinaddr[2]\ : SLE
      port map(D => \rbinaddr_3[2]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[2]_net_1\);
    
    \wsync1_rptr[31]\ : SLE
      port map(D => \raddr_gray[31]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[31]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[32]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIPD1S9_S[32]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[32]\);
    
    \wbinaddr_RNIJ33O8[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_28, S
         => \wbinaddr_RNIJ33O8_S[29]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_29);
    
    \wsync1_rptr[8]\ : SLE
      port map(D => \raddr_gray[8]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[8]_net_1\);
    
    \rbinaddr[18]\ : SLE
      port map(D => \rbinaddr_3[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[18]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_93\ : ARI1
      generic map(INIT => x"60609")

      port map(A => \rsync2_wptr[4]_net_1\, B => 
        \rbinaddr_RNI4EE41_S[4]\, C => \rbinaddr_RNII5581_S[5]\, 
        D => fifo_empty_xhdl3_0_N_6, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[1]\, S => OPEN, Y => OPEN, 
        FCO => \fifo_empty_xhdl3_0_data_tmp[2]\);
    
    \wbinaddr[16]\ : SLE
      port map(D => \wbinaddr_2[16]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[16]_net_1\);
    
    \Write_Bin_Ptr.wbinaddr_2[16]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIHJPS3_S[16]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[16]\);
    
    \waddr_gray[18]\ : SLE
      port map(D => \wgraynext[18]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[18]_net_1\);
    
    \rbinaddr_RNI03P48[29]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[29]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_28, S
         => \rbinaddr_RNI03P48_S[29]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_29);
    
    \rgraynext[21]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIPCKS5_S[22]\, B => 
        \rbinaddr_RNISMAI5_S[21]\, Y => \rgraynext[21]_net_1\);
    
    \wbinaddr[14]\ : SLE
      port map(D => \wbinaddr_2[14]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[14]_net_1\);
    
    \rbinaddr[11]\ : SLE
      port map(D => \rbinaddr_3[11]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rbinaddr[11]_net_1\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_46\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNIVVSU3_S[16]\, B => 
        \rsync2_wptr[15]_net_1\, C => \rbinaddr_RNIV7KK3_S[15]\, 
        Y => fifo_empty_xhdl3_0_N_46);
    
    \rgraynext[23]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNIMR7H6_S[24]\, B => 
        \rbinaddr_RNIN3U66_S[23]\, Y => \rgraynext[23]_net_1\);
    
    \rgraynext[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI2R203_S[13]\, B => 
        \rbinaddr_RNI56QL2_S[12]\, Y => \rgraynext[12]_net_1\);
    
    \rbinaddr_RNIKD0N1[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_8, S
         => \rbinaddr_RNIKD0N1_S[9]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_9);
    
    \Write_Bin_Ptr.wbinaddr_2[30]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNIKG249_S[30]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[30]\);
    
    \Read_Bin_Ptr.rbinaddr_3[19]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI5ENT4_S[19]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[19]\);
    
    \rbinaddr_RNI0EAP[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_0, S
         => \rbinaddr_RNI0EAP_S[1]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_1);
    
    \rsync1_wptr[12]\ : SLE
      port map(D => \waddr_gray[12]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rsync1_wptr[12]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[11]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI9IHB2_S[11]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[11]\);
    
    \raddr_gray[2]\ : SLE
      port map(D => \rgraynext[2]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \raddr_gray[2]_net_1\);
    
    \waddr_gray[20]\ : SLE
      port map(D => \wgraynext[20]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[20]_net_1\);
    
    \wgraynext[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNIM4P31_S[7]\, B => 
        \wbinaddr_RNI1PV01_S[6]\, Y => \wgraynext[6]_net_1\);
    
    \rgraynext[18]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rbinaddr_RNI5ENT4_S[19]\, B => 
        \rbinaddr_RNI2JEJ4_S[18]\, Y => \rgraynext[18]_net_1\);
    
    \rbinaddr_RNIEV812[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_9, S
         => \rbinaddr_RNIEV812_S[10]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_10);
    
    \wsync2_rptr[4]\ : SLE
      port map(D => \wsync1_rptr[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync2_rptr[4]_net_1\);
    
    \wgraynext[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI289L1_S[10]\, B => 
        \wbinaddr_RNI3VB91_S[9]\, Y => \wgraynext[9]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[10]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIEV812_S[10]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[10]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_16\ : CFG3
      generic map(INIT => x"96")

      port map(A => \rbinaddr_RNISO3F8_S[30]\, B => 
        \rsync2_wptr[29]_net_1\, C => \rbinaddr_RNI03P48_S[29]\, 
        Y => fifo_empty_xhdl3_0_N_71);
    
    \Write_Bin_Ptr.wbinaddr_2[6]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \wbinaddr_RNI1PV01_S[6]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \wbinaddr_2[6]\);
    
    \Read_Bin_Ptr.rbinaddr_3[27]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNIP95G7_S[27]\, B => hsel2_0_a2_1, 
        C => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[27]\);
    
    \Gen_Empty.fifo_empty_xhdl3_0_I_99\ : ARI1
      generic map(INIT => x"69900")

      port map(A => VCC_net_1, B => \rbinaddr_RNIN7P39_S[32]\, C
         => \rsync2_wptr[32]_net_1\, D => GND_net_1, FCI => 
        \fifo_empty_xhdl3_0_data_tmp[15]\, S => OPEN, Y => OPEN, 
        FCO => fifo_empty_xhdl3_0_N_2);
    
    \wbinaddr_RNI3T3D2[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_11, S
         => \wbinaddr_RNI3T3D2_S[12]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_12);
    
    \waddr_gray[15]\ : SLE
      port map(D => \wgraynext[15]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[15]_net_1\);
    
    \waddr_gray[0]\ : SLE
      port map(D => \wgraynext[0]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[0]_net_1\);
    
    \Read_Bin_Ptr.rbinaddr_3[1]\ : CFG4
      generic map(INIT => x"AA2A")

      port map(A => \rbinaddr_RNI0EAP_S[1]\, B => hsel2_0_a2_1, C
         => masterAddrInProg_0, D => valid_ahbcmd_i_o3_1, Y => 
        \rbinaddr_3[1]\);
    
    \rbinaddr_RNI0P594[17]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[17]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_16, S
         => \rbinaddr_RNI0P594_S[17]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_17);
    
    \wgraynext[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wbinaddr_RNI2I612_S[11]\, B => 
        \wbinaddr_RNI289L1_S[10]\, Y => \wgraynext[10]_net_1\);
    
    \wbinaddr_RNI67I05[19]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wbinaddr[19]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_wbinnext_cry_18, S
         => \wbinaddr_RNI67I05_S[19]\, Y => OPEN, FCO => 
        un3_wbinnext_cry_19);
    
    \wbinaddr[0]\ : SLE
      port map(D => \wbinaddr_2[0]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wbinaddr[0]_net_1\);
    
    \waddr_gray[3]\ : SLE
      port map(D => \wgraynext[3]_net_1\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[3]_net_1\);
    
    \rbinaddr_RNIHNIF1[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rbinaddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => un3_rbinnext_cry_6, S
         => \rbinaddr_RNIHNIF1_S[7]\, Y => OPEN, FCO => 
        un3_rbinnext_cry_7);
    
    \waddr_gray[26]\ : SLE
      port map(D => \wgraynext[26]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \waddr_gray[26]_net_1\);
    
    \wsync1_rptr[32]\ : SLE
      port map(D => \raddr_gray[32]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wsync1_rptr[32]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Synchronizer_AXItoAHBHX is

    port( synchronizer_1_0                   : out   std_logic;
          BVALID_sync                        : out   std_logic;
          axi_read_rlast                     : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID : in    std_logic;
          post_sync_1_reg                    : out   std_logic;
          SDRCLK_c                           : in    std_logic;
          ARESET_n                           : in    std_logic
        );

end Synchronizer_AXItoAHBHX;

architecture DEF_ARCH of Synchronizer_AXItoAHBHX is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \pre_sync_0_reg\, VCC_net_1, \pre_sync_0_reg_0\, 
        GND_net_1, \synchronizer_0[0]_net_1\, 
        \synchronizer_0[1]_net_1\, \synchronizer_1_0\, 
        \synchronizer_1[1]_net_1\, \pre_sync_1_reg\, 
        \post_sync_0_reg\, \pre_sync_1_reg_0\ : std_logic;

begin 

    synchronizer_1_0 <= \synchronizer_1_0\;

    \synchronizer_1[1]\ : SLE
      port map(D => \pre_sync_1_reg\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_1[1]_net_1\);
    
    pre_sync_0_reg : SLE
      port map(D => \pre_sync_0_reg_0\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pre_sync_0_reg\);
    
    \synchronizer_0[1]\ : SLE
      port map(D => \pre_sync_0_reg\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_0[1]_net_1\);
    
    pre_sync_1_reg : SLE
      port map(D => \pre_sync_1_reg_0\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \pre_sync_1_reg\);
    
    pre_sync_0_reg_0 : CFG2
      generic map(INIT => x"6")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_BVALID, B => 
        \pre_sync_0_reg\, Y => \pre_sync_0_reg_0\);
    
    \synchronizer_1[0]\ : SLE
      port map(D => \synchronizer_1[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_1_0\);
    
    \synchronizer_0[0]\ : SLE
      port map(D => \synchronizer_0[1]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \synchronizer_0[0]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    post_sync_0_reg : SLE
      port map(D => \synchronizer_0[0]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \post_sync_0_reg\);
    
    Dout_0 : CFG2
      generic map(INIT => x"6")

      port map(A => \synchronizer_0[0]_net_1\, B => 
        \post_sync_0_reg\, Y => BVALID_sync);
    
    pre_sync_1_reg_0 : CFG2
      generic map(INIT => x"6")

      port map(A => \pre_sync_1_reg\, B => axi_read_rlast, Y => 
        \pre_sync_1_reg_0\);
    
    \post_sync_1_reg\ : SLE
      port map(D => \synchronizer_1_0\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        post_sync_1_reg);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_AXIAccessControlHX is

    port( COREAHBLTOAXI_0_AXIMasterIF_WDATA    : out   std_logic_vector(63 downto 16);
          rdch_fifo_wr_data                    : out   std_logic_vector(31 downto 0);
          HADDR_d                              : in    std_logic_vector(27 downto 0);
          HSIZE_d                              : in    std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : in    std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : out   std_logic_vector(27 downto 1);
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : out   std_logic_vector(1 downto 0);
          axi_current_state_0                  : out   std_logic;
          axi_current_state_3                  : out   std_logic;
          axi_current_state_2                  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : out   std_logic;
          N_1448_i                             : out   std_logic;
          N_1449_i                             : out   std_logic;
          N_1450_i                             : out   std_logic;
          N_202_i                              : out   std_logic;
          N_201_i                              : out   std_logic;
          N_200_i                              : out   std_logic;
          N_197_i                              : out   std_logic;
          N_195_i                              : out   std_logic;
          N_134_i                              : out   std_logic;
          N_133_i                              : out   std_logic;
          N_380_i                              : out   std_logic;
          N_278_i                              : out   std_logic;
          N_381_i                              : out   std_logic;
          N_382_i                              : out   std_logic;
          N_277_i                              : out   std_logic;
          N_276_i                              : out   std_logic;
          N_275_i                              : out   std_logic;
          N_274_i                              : out   std_logic;
          N_273_i                              : out   std_logic;
          N_272_i                              : out   std_logic;
          N_203_i                              : out   std_logic;
          N_137_i                              : out   std_logic;
          N_136_i                              : out   std_logic;
          N_135_i                              : out   std_logic;
          N_209                                : in    std_logic;
          N_217                                : in    std_logic;
          N_210                                : in    std_logic;
          N_218                                : in    std_logic;
          N_213                                : in    std_logic;
          N_221                                : in    std_logic;
          N_214                                : in    std_logic;
          N_222                                : in    std_logic;
          N_215                                : in    std_logic;
          N_223                                : in    std_logic;
          N_432                                : in    std_logic;
          N_439                                : in    std_logic;
          N_431                                : in    std_logic;
          N_438                                : in    std_logic;
          N_430                                : in    std_logic;
          N_437                                : in    std_logic;
          N_429                                : in    std_logic;
          N_436                                : in    std_logic;
          N_428                                : in    std_logic;
          N_435                                : in    std_logic;
          N_427                                : in    std_logic;
          N_434                                : in    std_logic;
          N_426                                : in    std_logic;
          N_433                                : in    std_logic;
          N_421                                : in    std_logic;
          N_425                                : in    std_logic;
          N_420                                : in    std_logic;
          N_424                                : in    std_logic;
          N_419                                : in    std_logic;
          N_423                                : in    std_logic;
          N_418                                : in    std_logic;
          N_422                                : in    std_logic;
          N_417                                : in    std_logic;
          N_414                                : in    std_logic;
          N_416                                : in    std_logic;
          N_413                                : in    std_logic;
          N_328                                : in    std_logic;
          N_440                                : in    std_logic;
          N_412                                : in    std_logic;
          N_415                                : in    std_logic;
          N_410                                : in    std_logic;
          N_411                                : in    std_logic;
          N_286                                : in    std_logic;
          N_293                                : in    std_logic;
          N_285                                : in    std_logic;
          N_292                                : in    std_logic;
          N_284                                : in    std_logic;
          N_291                                : in    std_logic;
          N_283                                : in    std_logic;
          N_290                                : in    std_logic;
          N_282                                : in    std_logic;
          N_289                                : in    std_logic;
          N_281                                : in    std_logic;
          N_288                                : in    std_logic;
          N_151                                : in    std_logic;
          N_160                                : in    std_logic;
          N_150                                : in    std_logic;
          N_159                                : in    std_logic;
          N_149                                : in    std_logic;
          N_158                                : in    std_logic;
          N_148                                : in    std_logic;
          N_157                                : in    std_logic;
          N_147                                : in    std_logic;
          N_156                                : in    std_logic;
          N_1451_i                             : out   std_logic;
          N_1447_i                             : out   std_logic;
          N_1452_i                             : out   std_logic;
          N_1446_i                             : out   std_logic;
          wready_m_xhdl2                       : in    std_logic;
          N_73_i_0                             : out   std_logic;
          N_72_i                               : out   std_logic;
          N_1445_i                             : out   std_logic;
          N_48                                 : out   std_logic;
          N_75_i                               : out   std_logic;
          ahb_wr_done_sync                     : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic;
          N_98                                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : in    std_logic;
          araddr_arvalid_clr_d                 : out   std_logic;
          awaddr_awvalid_clr_d                 : out   std_logic;
          ahb_rd_req_sync                      : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : in    std_logic;
          latch_ahb_sig_sync                   : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : out   std_logic;
          rdch_fifo_wr_en_r                    : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : out   std_logic;
          axi_read_rlast                       : out   std_logic;
          HMASTLOCK_d                          : in    std_logic;
          HWRITE_d                             : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          ARESET_n                             : in    std_logic
        );

end CoreAHBLtoAXI_AXIAccessControlHX;

architecture DEF_ARCH of CoreAHBLtoAXI_AXIAccessControlHX is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \swap_rd_data_byte[2]_net_1\, VCC_net_1, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, GND_net_1, 
        \AWADDR_incr[0]_net_1\, \AWADDR_incr_9_i_m2[0]_net_1\, 
        \AWADDR_incr[1]_net_1\, \AWADDR_incr_9_i_m2[1]_net_1\, 
        \AWADDR_incr[2]_net_1\, \AWADDR_incr_9_i_m2[2]_net_1\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, \HSIZE_sync_150\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, \HSIZE_sync_151\, 
        \burstcount_reg[0]_net_1\, N_93_i, 
        \burstcount_reg[1]_net_1\, N_68_i, 
        \burstcount_reg[2]_net_1\, N_69_i, 
        \burstcount_reg[3]_net_1\, \SUM_i_m3[3]\, 
        \burstcount_reg[4]_net_1\, N_70_i_0, \store_ahb_sig\, 
        \rdch_write_data_r[63]_net_1\, 
        \axi_read_data_xhdl68_1_i_i_a3\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, \HADDR_sync_153\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, \HADDR_sync_154\, 
        \HADDR_sync_155\, \rdch_write_data_r[48]_net_1\, 
        \rdch_write_data_r[49]_net_1\, 
        \rdch_write_data_r[50]_net_1\, 
        \rdch_write_data_r[51]_net_1\, 
        \rdch_write_data_r[52]_net_1\, 
        \rdch_write_data_r[53]_net_1\, 
        \rdch_write_data_r[54]_net_1\, 
        \rdch_write_data_r[55]_net_1\, 
        \rdch_write_data_r[56]_net_1\, 
        \rdch_write_data_r[57]_net_1\, 
        \rdch_write_data_r[58]_net_1\, 
        \rdch_write_data_r[59]_net_1\, 
        \rdch_write_data_r[60]_net_1\, 
        \rdch_write_data_r[61]_net_1\, 
        \rdch_write_data_r[62]_net_1\, 
        \rdch_write_data_r[33]_net_1\, 
        \rdch_write_data_r[34]_net_1\, 
        \rdch_write_data_r[35]_net_1\, 
        \rdch_write_data_r[36]_net_1\, 
        \rdch_write_data_r[37]_net_1\, 
        \rdch_write_data_r[38]_net_1\, 
        \rdch_write_data_r[39]_net_1\, 
        \rdch_write_data_r[40]_net_1\, 
        \rdch_write_data_r[41]_net_1\, 
        \rdch_write_data_r[42]_net_1\, 
        \rdch_write_data_r[43]_net_1\, 
        \rdch_write_data_r[44]_net_1\, 
        \rdch_write_data_r[45]_net_1\, 
        \rdch_write_data_r[46]_net_1\, 
        \rdch_write_data_r[47]_net_1\, 
        \rdch_write_data_r[18]_net_1\, 
        \rdch_write_data_r[19]_net_1\, 
        \rdch_write_data_r[20]_net_1\, 
        \rdch_write_data_r[21]_net_1\, 
        \rdch_write_data_r[22]_net_1\, 
        \rdch_write_data_r[23]_net_1\, 
        \rdch_write_data_r[24]_net_1\, 
        \rdch_write_data_r[25]_net_1\, 
        \rdch_write_data_r[26]_net_1\, 
        \rdch_write_data_r[27]_net_1\, 
        \rdch_write_data_r[28]_net_1\, 
        \rdch_write_data_r[29]_net_1\, 
        \rdch_write_data_r[30]_net_1\, 
        \rdch_write_data_r[31]_net_1\, 
        \rdch_write_data_r[32]_net_1\, 
        \rdch_write_data_r[3]_net_1\, 
        \rdch_write_data_r[4]_net_1\, 
        \rdch_write_data_r[5]_net_1\, 
        \rdch_write_data_r[6]_net_1\, 
        \rdch_write_data_r[7]_net_1\, 
        \rdch_write_data_r[8]_net_1\, 
        \rdch_write_data_r[9]_net_1\, 
        \rdch_write_data_r[10]_net_1\, 
        \rdch_write_data_r[11]_net_1\, 
        \rdch_write_data_r[12]_net_1\, 
        \rdch_write_data_r[13]_net_1\, 
        \rdch_write_data_r[14]_net_1\, 
        \rdch_write_data_r[15]_net_1\, 
        \rdch_write_data_r[16]_net_1\, 
        \rdch_write_data_r[17]_net_1\, 
        \rdch_write_data_r[0]_net_1\, 
        \rdch_write_data_r[1]_net_1\, 
        \rdch_write_data_r[2]_net_1\, \wvalid_reg\, N_99_i, 
        \wvalid_reg_1_sqmuxa_i_0\, \HWRITE_sync\, 
        \axi_wstrb[9]_net_1\, N_1737_i, \axi_wstrb[8]_net_1\, 
        N_1739_i, \axi_wstrb[7]_net_1\, N_1741_i, 
        \axi_wstrb[6]_net_1\, \axi_wstrb_ns_i_i[19]_net_1\, 
        \axi_wstrb[5]_net_1\, N_1745_i, \axi_wstrb[4]_net_1\, 
        N_1747_i, \axi_wstrb[3]_net_1\, N_1749_i, 
        \axi_wstrb[2]_net_1\, N_1751_i, \axi_wstrb[1]_net_1\, 
        N_1753_i, \axi_wstrb[0]_net_1\, N_1755_i, 
        \axi_wstrb[24]_net_1\, N_1708_i, \axi_wstrb[23]_net_1\, 
        N_1710_i, \axi_wstrb[22]_net_1\, N_383_i, 
        \axi_wstrb[21]_net_1\, N_1713_i, \axi_wstrb[20]_net_1\, 
        N_1715_i, \axi_wstrb[19]_net_1\, N_1717_i, 
        \axi_wstrb[18]_net_1\, N_1719_i, \axi_wstrb[17]_net_1\, 
        N_1721_i, \axi_wstrb[16]_net_1\, N_1723_i, 
        \axi_wstrb[15]_net_1\, N_1725_i, \axi_wstrb[14]_net_1\, 
        N_1727_i, \axi_wstrb[13]_net_1\, N_1729_i, 
        \axi_wstrb[12]_net_1\, N_1731_i, \axi_wstrb[11]_net_1\, 
        N_1733_i, \axi_wstrb[10]_net_1\, N_1735_i, 
        \axi_current_state[2]_net_1\, \axi_current_state_ns[3]\, 
        \axi_current_state_0\, \axi_current_state_ns[4]\, 
        \axi_current_state[0]_net_1\, \axi_current_state_ns[5]\, 
        \axi_current_state[5]_net_1\, \axi_current_state_ns[0]\, 
        \axi_current_state_3\, \axi_current_state_ns[1]\, 
        \axi_current_state_2\, \axi_current_state_ns[2]\, 
        \wvalid_set_r\, wvalid_set_r_1, axi_read_rlast_xhdl26_1, 
        \COREAHBLTOAXI_0_AXIMasterIF_RREADY\, 
        \rready_set_xhdl69_1_i_i\, \wvalid_clr_t\, WLAST, 
        \COREAHBLTOAXI_0_AXIMasterIF_WVALID\, temp_xhdl42, 
        \latch_ahb_sig_sync_d\, \wvalid_reg_r\, \BVALID_reg\, 
        \ahb_rd_req_sync_d\, awaddr_awvalid_clr_d_net_1, N_88_i, 
        araddr_arvalid_clr_d_net_1, N_274_i_0, N_279, N_265, 
        N_280, N_552, N_71_i_1, 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_1_i_0\, N_71_i, 
        \un1_axi_current_state_5_i_o3_sx\, N_82, N_396, 
        \WDATA_i_i_o2_1[25]_net_1\, N_390, N_551, 
        \WDATA_i_o2_i_m2_1[31]_net_1\, N_330, N_48_i, 
        \un34_i_a2_4_a2_0[2]_net_1\, N_558, N_271, N_397, N_83, 
        N_79, latch_wr_resp_set_xhdl66_0_sqmuxa, N_555, N_395, 
        N_394, N_100_i, un1_axi_current_state_i, 
        \un34_i_a2_5_a2_2[3]_net_1\, \un34_i_a2_5_a2_1[4]_net_1\, 
        \un34_i_a2_0_a2_1[1]_net_1\, 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_i_0\, 
        \un34_i_a2_5_a2_2[5]_net_1\, \un34_i_a2_4_a2_2[6]_net_1\, 
        N_105, N_115, N_550, N_67_i_0, N_91, N_81, N_523_1, 
        \axi_wstrb_ns_i_0_0[15]_net_1\, N_442, N_443, N_445, 
        N_446, N_444, N_441, \SUM_i_o3_0[4]\, 
        \axi_wstrb_ns_i_0_0[6]_net_1\, 
        \axi_wstrb_ns_i_0_0[18]_net_1\, N_194, N_373, N_388, 
        N_389, N_1723_1, N_86, N_140, 
        \un1_rd_data_c_xhdl44_1_sqmuxa_i_0\, \N_72_i\, N_392, 
        N_346, N_384, WDATA_sn_N_17_mux, N_563, N_139, N_142
         : std_logic;

begin 

    COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2) <= 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\;
    COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1) <= 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\;
    COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1) <= 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\;
    COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0) <= 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\;
    axi_current_state_0 <= \axi_current_state_0\;
    axi_current_state_3 <= \axi_current_state_3\;
    axi_current_state_2 <= \axi_current_state_2\;
    N_72_i <= \N_72_i\;
    araddr_arvalid_clr_d <= araddr_arvalid_clr_d_net_1;
    awaddr_awvalid_clr_d <= awaddr_awvalid_clr_d_net_1;
    COREAHBLTOAXI_0_AXIMasterIF_WVALID <= 
        \COREAHBLTOAXI_0_AXIMasterIF_WVALID\;
    COREAHBLTOAXI_0_AXIMasterIF_RREADY <= 
        \COREAHBLTOAXI_0_AXIMasterIF_RREADY\;

    \WDATA_0[29]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_432, B => N_439, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(29));
    
    \HADDR_sync[11]\ : SLE
      port map(D => HADDR_d(11), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11));
    
    \axi_wstrb_RNO[21]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => N_441, C => N_395, Y => N_1713_i);
    
    \WDATA_i_o4_i_o2_RNI7PUD3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_283, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_290, Y => N_274_i);
    
    \WDATA_0[44]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_290, B => N_194, C => N_142, D => N_283, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(44));
    
    \axi_wstrb_RNO[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[3]_net_1\, Y => 
        N_1749_i);
    
    \WDATA_0_0[47]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_415, B => N_194, C => N_142, D => N_412, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(47));
    
    \rdch_write_data_r[1]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(1), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[1]_net_1\);
    
    \rdch_fifo_wr_data[27]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[59]_net_1\, B => 
        \rdch_write_data_r[27]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(27));
    
    wvalid_set_r : SLE
      port map(D => wvalid_set_r_1, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wvalid_set_r\);
    
    \burstcount_reg[4]\ : SLE
      port map(D => N_70_i_0, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \burstcount_reg[4]_net_1\);
    
    \WDATA_1[61]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_439, B => N_140, C => N_139, D => N_432, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(61));
    
    \burstcount_reg[0]\ : SLE
      port map(D => N_93_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \burstcount_reg[0]_net_1\);
    
    \axi_wstrb_ns_i_0_o2[6]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, Y => N_271);
    
    \WDATA_i_o2_i[31]\ : CFG3
      generic map(INIT => x"F9")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_330, 
        Y => N_373);
    
    \WDATA_0_o2_0_o2_0_RNI9QGA1[36]\ : CFG3
      generic map(INIT => x"A2")

      port map(A => N_551, B => N_397, C => N_388, Y => 
        WDATA_sn_N_17_mux);
    
    \un34_i_a2_4_a2_0_0_RNIEMD41[2]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \axi_wstrb[12]_net_1\, B => 
        \un34_i_a2_4_a2_0[2]_net_1\, C => N_558, D => N_563, Y
         => N_1450_i);
    
    \WDATA_i_o4_i_o2_RNI3LUD3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_285, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_292, Y => N_276_i);
    
    \axi_wstrb_ns_i_0_m2[12]\ : CFG4
      generic map(INIT => x"F044")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, C => 
        \axi_wstrb[13]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_445);
    
    \axi_wstrb_RNO[12]\ : CFG4
      generic map(INIT => x"0604")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_446, 
        D => N_395, Y => N_1731_i);
    
    HADDR_sync_155 : CFG4
      generic map(INIT => x"E4F0")

      port map(A => \latch_ahb_sig_sync_d\, B => HADDR_d(2), C
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, D => 
        latch_ahb_sig_sync, Y => \HADDR_sync_155\);
    
    \axi_wstrb[11]\ : SLE
      port map(D => N_1733_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[11]_net_1\);
    
    \axi_wstrb_RNO[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[8]_net_1\, Y => 
        N_1739_i);
    
    \rdch_write_data_r[6]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(6), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[6]_net_1\);
    
    \axi_wstrb_RNO[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[9]_net_1\, Y => 
        N_1737_i);
    
    \axi_wstrb[8]\ : SLE
      port map(D => N_1739_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[8]_net_1\);
    
    wvalid_reg_r : SLE
      port map(D => \wvalid_reg\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wvalid_reg_r\);
    
    \un34_i_a2_0_a2_0[0]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \axi_wstrb[3]_net_1\, B => 
        \axi_wstrb[2]_net_1\, C => \axi_wstrb[1]_net_1\, D => 
        \axi_wstrb[0]_net_1\, Y => N_552);
    
    \rdch_fifo_wr_data[23]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[55]_net_1\, B => 
        \rdch_write_data_r[23]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(23));
    
    \axi_wstrb_RNO[17]\ : CFG4
      generic map(INIT => x"0A03")

      port map(A => \axi_wstrb[17]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, C => N_394, D
         => N_395, Y => N_1721_i);
    
    \axi_wstrb[21]\ : SLE
      port map(D => N_1713_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[21]_net_1\);
    
    \WDATA_i_o4_i_o2_RNIDVUD3[4]\ : CFG4
      generic map(INIT => x"00D8")

      port map(A => N_396, B => N_415, C => N_412, D => 
        WDATA_sn_N_17_mux, Y => N_203_i);
    
    \axi_current_state_ns_0[4]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARREADY, B => 
        N_115, C => \axi_current_state_0\, Y => 
        \axi_current_state_ns[4]\);
    
    \HADDR_sync[18]\ : SLE
      port map(D => HADDR_d(18), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18));
    
    \AWADDR_incr_9_i_m2[0]\ : CFG4
      generic map(INIT => x"AAC3")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, B
         => \AWADDR_incr[0]_net_1\, C => N_279, D => N_48_i, Y
         => \AWADDR_incr_9_i_m2[0]_net_1\);
    
    \un34_i_a2_5_a2_0_RNI1F3H[5]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => N_550, B => \un34_i_a2_5_a2_2[5]_net_1\, C
         => \axi_wstrb[17]_net_1\, D => \axi_wstrb[14]_net_1\, Y
         => N_1447_i);
    
    \rdch_write_data_r[38]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(38), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[38]_net_1\);
    
    \un1_burstcount_reg_2_1.SUM_i_m3[3]\ : CFG3
      generic map(INIT => x"09")

      port map(A => N_86, B => \burstcount_reg[3]_net_1\, C => 
        N_79, Y => \SUM_i_m3[3]\);
    
    \rdch_fifo_wr_data[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[34]_net_1\, B => 
        \rdch_write_data_r[2]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(2));
    
    \rdch_fifo_wr_data[21]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[53]_net_1\, B => 
        \rdch_write_data_r[21]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(21));
    
    wvalid_reg_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"8F88")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_WREADY, B => 
        WLAST, C => \wvalid_clr_t\, D => \axi_current_state_2\, Y
         => \wvalid_reg_1_sqmuxa_i_0\);
    
    rdch_fifo_wr_en_r_xhdl24 : SLE
      port map(D => \axi_read_data_xhdl68_1_i_i_a3\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rdch_fifo_wr_en_r);
    
    \rdch_write_data_r[31]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(31), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[31]_net_1\);
    
    \axi_wstrb_RNO[13]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => N_445, C => N_395, Y => N_1729_i);
    
    \un1_burstcount_reg_2_1.SUM_i_o3[2]\ : CFG3
      generic map(INIT => x"FB")

      port map(A => \burstcount_reg[0]_net_1\, B => N_67_i_0, C
         => \burstcount_reg[1]_net_1\, Y => N_91);
    
    \axi_current_state_ns_0[1]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_AWREADY, B => 
        \axi_current_state_3\, C => ahb_wr_done_sync, D => 
        \axi_current_state[5]_net_1\, Y => 
        \axi_current_state_ns[1]\);
    
    \un1_burstcount_reg_2_1.SUM_i_o3_0[4]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \burstcount_reg[3]_net_1\, B => 
        \burstcount_reg[2]_net_1\, C => \burstcount_reg[1]_net_1\, 
        D => \burstcount_reg[0]_net_1\, Y => \SUM_i_o3_0[4]\);
    
    \WDATA_i_o4_i_o2_RNIVJJK3[4]\ : CFG4
      generic map(INIT => x"00D8")

      port map(A => N_396, B => N_434, C => N_427, D => 
        WDATA_sn_N_17_mux, Y => N_381_i);
    
    \rdch_write_data_r[49]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(49), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[49]_net_1\);
    
    \axi_wstrb_ns_i_0_o2[8]\ : CFG2
      generic map(INIT => x"B")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_394);
    
    \WDATA_i_o4_i_o2_RNI5NUD3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_284, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_291, Y => N_275_i);
    
    \WDATA_i_o2_i_RNIPFPG3[31]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_217, B => N_209, C => WDATA_sn_N_17_mux, D
         => N_373, Y => N_195_i);
    
    \axi_wstrb_ns_i_0_m2[7]\ : CFG3
      generic map(INIT => x"8D")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => N_271, C => \axi_wstrb[18]_net_1\, Y => N_442);
    
    \axi_wstrb_RNO[20]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[20]_net_1\, Y => 
        N_1715_i);
    
    wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"777F")

      port map(A => \wvalid_set_r\, B => \wvalid_reg\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_i_0\);
    
    \axi_wstrb_RNO[18]\ : CFG4
      generic map(INIT => x"0600")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, C => N_442, 
        D => N_395, Y => N_1719_i);
    
    \axi_wstrb[4]\ : SLE
      port map(D => N_1747_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[4]_net_1\);
    
    \HADDR_sync[20]\ : SLE
      port map(D => HADDR_d(20), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20));
    
    \axi_current_state[3]\ : SLE
      port map(D => \axi_current_state_ns[2]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state_2\);
    
    \rdch_write_data_r[23]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(23), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[23]_net_1\);
    
    \WDATA_1_0[62]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_440, B => N_140, C => N_139, D => N_328, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(62));
    
    \rdch_write_data_r[50]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(50), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[50]_net_1\);
    
    \axi_wstrb[9]\ : SLE
      port map(D => N_1737_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[9]_net_1\);
    
    \un1_burstcount_reg_2_1.N_70_i\ : CFG4
      generic map(INIT => x"2122")

      port map(A => \burstcount_reg[4]_net_1\, B => N_79, C => 
        \SUM_i_o3_0[4]\, D => N_67_i_0, Y => N_70_i_0);
    
    \axi_current_state_ns_0[3]\ : CFG4
      generic map(INIT => x"2F22")

      port map(A => \axi_current_state_2\, B => N_82, C => 
        \BVALID_reg\, D => \axi_current_state[2]_net_1\, Y => 
        \axi_current_state_ns[3]\);
    
    \WDATA_i_o4_i_o2[4]\ : CFG2
      generic map(INIT => x"B")

      port map(A => N_394, B => \AWADDR_incr[2]_net_1\, Y => 
        N_396);
    
    BVALID_reg : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_BVALID, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \BVALID_reg\);
    
    \axi_wstrb[15]\ : SLE
      port map(D => N_1725_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[15]_net_1\);
    
    \un1_burstcount_reg_2_1.SUM_i_o3[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \axi_current_state_3\, B => 
        \axi_current_state_0\, Y => N_79);
    
    \WDATA_0[39]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_434, B => N_194, C => N_142, D => N_427, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(39));
    
    \rdch_write_data_r[10]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(10), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[10]_net_1\);
    
    \axi_current_state[2]\ : SLE
      port map(D => \axi_current_state_ns[3]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state[2]_net_1\);
    
    \WDATA_1[54]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_436, B => N_140, C => N_139, D => N_429, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(54));
    
    temp_xhdl42_0 : CFG4
      generic map(INIT => x"22A2")

      port map(A => \wvalid_reg\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, C => 
        \axi_current_state_ns[2]\, D => WLAST, Y => temp_xhdl42);
    
    \rdch_write_data_r[24]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(24), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[24]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \axi_wstrb[3]\ : SLE
      port map(D => N_1749_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[3]_net_1\);
    
    \rdch_fifo_wr_data[24]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[56]_net_1\, B => 
        \rdch_write_data_r[24]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(24));
    
    \rdch_write_data_r[27]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(27), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[27]_net_1\);
    
    wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_1_i_0 : CFG4
      generic map(INIT => x"FFF7")

      port map(A => \wvalid_set_r\, B => \wvalid_reg\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_1_i_0\);
    
    \rdch_write_data_r[61]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(61), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[61]_net_1\);
    
    \axi_wstrb[12]\ : SLE
      port map(D => N_1731_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[12]_net_1\);
    
    \AWADDR_incr_9_i_m2[2]\ : CFG4
      generic map(INIT => x"AAC3")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \AWADDR_incr[2]_net_1\, C => N_346, D => N_48_i, Y
         => \AWADDR_incr_9_i_m2[2]_net_1\);
    
    \rdch_fifo_wr_data[16]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[48]_net_1\, B => 
        \rdch_write_data_r[16]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(16));
    
    \HADDR_sync[3]\ : SLE
      port map(D => HADDR_d(3), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3));
    
    \axi_current_state_ns_0[5]\ : CFG4
      generic map(INIT => x"BA30")

      port map(A => \axi_current_state[0]_net_1\, B => 
        \HWRITE_sync\, C => N_81, D => N_83, Y => 
        \axi_current_state_ns[5]\);
    
    un1_rd_data_c_xhdl44_1_sqmuxa_i_0 : CFG4
      generic map(INIT => x"AF11")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \swap_rd_data_byte[2]_net_1\, C => N_555, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => 
        \un1_rd_data_c_xhdl44_1_sqmuxa_i_0\);
    
    \rdch_write_data_r[52]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(52), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[52]_net_1\);
    
    \rdch_fifo_wr_data[19]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[51]_net_1\, B => 
        \rdch_write_data_r[19]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(19));
    
    \HADDR_sync[4]\ : SLE
      port map(D => HADDR_d(4), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4));
    
    \WDATA_1[60]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_218, B => N_140, C => N_139, D => N_210, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(60));
    
    \axi_current_state_ns_0_a3_0[4]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \axi_current_state[5]_net_1\, B => 
        ahb_rd_req_sync, C => \ahb_rd_req_sync_d\, D => 
        ahb_wr_done_sync, Y => N_115);
    
    un1_axi_current_state_i_0_a2_0_a3 : CFG3
      generic map(INIT => x"01")

      port map(A => \axi_current_state_3\, B => 
        \axi_current_state[2]_net_1\, C => 
        \axi_current_state[5]_net_1\, Y => 
        un1_axi_current_state_i);
    
    \HADDR_sync[10]\ : SLE
      port map(D => HADDR_d(10), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10));
    
    \HADDR_sync[23]\ : SLE
      port map(D => HADDR_d(23), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23));
    
    \axi_wstrb[22]\ : SLE
      port map(D => N_383_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[22]_net_1\);
    
    \rdch_write_data_r[12]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(12), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[12]_net_1\);
    
    WVALID_xhdl11 : SLE
      port map(D => temp_xhdl42, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_WVALID\);
    
    \un1_burstcount_reg_2_1.N_93_i\ : CFG3
      generic map(INIT => x"BE")

      port map(A => N_79, B => N_67_i_0, C => 
        \burstcount_reg[0]_net_1\, Y => N_93_i);
    
    \HADDR_sync[0]\ : SLE
      port map(D => \HADDR_sync_153\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\);
    
    \axi_current_state_RNIGQJQ[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_ARREADY, B => 
        \axi_current_state_0\, Y => N_274_i_0);
    
    \rdch_write_data_r[39]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(39), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[39]_net_1\);
    
    un43_hburst_sync_i : CFG3
      generic map(INIT => x"DF")

      port map(A => \axi_current_state_3\, B => 
        awaddr_awvalid_clr_d_net_1, C => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, Y => N_48);
    
    \HADDR_sync[1]\ : SLE
      port map(D => \HADDR_sync_154\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\);
    
    \WDATA_i_o4_i_o2_RNIJ7JK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_150, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_159, Y => N_136_i);
    
    \WDATA_i_i_o2_1[25]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_551, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, Y => 
        \WDATA_i_i_o2_1[25]_net_1\);
    
    \WDATA_i_i_o2_0[25]\ : CFG3
      generic map(INIT => x"F1")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_194, 
        Y => N_392);
    
    \WDATA_0_a4_0_o2[36]\ : CFG4
      generic map(INIT => x"AF33")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \AWADDR_incr[2]_net_1\, C => N_271, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_194);
    
    \axi_wstrb_RNO[22]\ : CFG4
      generic map(INIT => x"0508")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \axi_wstrb[22]_net_1\, C => N_444, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_383_i);
    
    \axi_wstrb_ns_i_0_m2[4]\ : CFG4
      generic map(INIT => x"CC05")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, B
         => \axi_wstrb[21]_net_1\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_441);
    
    \WDATA_0_o2_0_o2[36]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => N_551, B => N_388, C => N_140, Y => N_142);
    
    \burstcount_reg_RNIPNJF[2]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \burstcount_reg[2]_net_1\, B => 
        \burstcount_reg[1]_net_1\, C => \burstcount_reg[0]_net_1\, 
        Y => N_71_i_1);
    
    \WDATA_0[23]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_430, B => N_437, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(23));
    
    \HADDR_sync[27]\ : SLE
      port map(D => HADDR_d(27), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27));
    
    \axi_wstrb_ns_i_0_0[6]\ : CFG4
      generic map(INIT => x"4E5F")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => N_271, C => \axi_wstrb[19]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, Y => 
        \axi_wstrb_ns_i_0_0[6]_net_1\);
    
    \axi_current_state_ns_0_a3[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \axi_current_state[2]_net_1\, B => 
        \BVALID_reg\, Y => latch_wr_resp_set_xhdl66_0_sqmuxa);
    
    \HADDR_sync[9]\ : SLE
      port map(D => HADDR_d(9), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9));
    
    \axi_wstrb[10]\ : SLE
      port map(D => N_1735_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[10]_net_1\);
    
    \HADDR_sync[22]\ : SLE
      port map(D => HADDR_d(22), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22));
    
    RREADY_xhdl20 : SLE
      port map(D => \rready_set_xhdl69_1_i_i\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_RREADY\);
    
    \WDATA_i_i[17]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_419, B => N_423, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(17));
    
    \axi_wstrb_RNO[7]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \axi_wstrb_ns_i_0_0[18]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_395, Y
         => N_1741_i);
    
    \axi_wstrb_RNIUBS7[24]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \axi_wstrb[24]_net_1\, B => 
        \axi_wstrb[22]_net_1\, C => \axi_wstrb[17]_net_1\, D => 
        \axi_wstrb[0]_net_1\, Y => N_1445_i);
    
    \HSIZE_sync_RNINK8N[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_551);
    
    \HADDR_sync[13]\ : SLE
      port map(D => HADDR_d(13), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13));
    
    \rdch_write_data_r[40]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(40), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[40]_net_1\);
    
    \axi_wstrb[2]\ : SLE
      port map(D => N_1751_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[2]_net_1\);
    
    \axi_wstrb[20]\ : SLE
      port map(D => N_1715_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[20]_net_1\);
    
    \AWADDR_incr_9_i_o2[0]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_WVALID\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_279);
    
    \WDATA_0_o2_0_o2_0[36]\ : CFG3
      generic map(INIT => x"A1")

      port map(A => \burstcount_reg[0]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, Y => N_388);
    
    \WDATA_i_o4_i_o2_RNIH5JK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_151, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_160, Y => N_137_i);
    
    \rdch_fifo_wr_data[6]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[38]_net_1\, B => 
        \rdch_write_data_r[6]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(6));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \rdch_write_data_r[3]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(3), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[3]_net_1\);
    
    \rdch_write_data_r[8]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(8), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[8]_net_1\);
    
    \axi_current_state[1]\ : SLE
      port map(D => \axi_current_state_ns[4]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state_0\);
    
    \axi_wstrb_RNO[23]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => N_443, C => N_395, Y => N_1710_i);
    
    \axi_wstrb[6]\ : SLE
      port map(D => \axi_wstrb_ns_i_i[19]_net_1\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[6]_net_1\);
    
    \rdch_fifo_wr_data[7]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[39]_net_1\, B => 
        \rdch_write_data_r[7]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(7));
    
    ARVALID : CFG2
      generic map(INIT => x"2")

      port map(A => \axi_current_state_0\, B => 
        araddr_arvalid_clr_d_net_1, Y => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID);
    
    \rdch_fifo_wr_data[8]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[40]_net_1\, B => 
        \rdch_write_data_r[8]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(8));
    
    \HADDR_sync[17]\ : SLE
      port map(D => HADDR_d(17), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17));
    
    \WDATA_1_0[57]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_416, B => N_140, C => N_139, D => N_413, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(57));
    
    \WDATA_1[59]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_438, B => N_140, C => N_139, D => N_431, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(59));
    
    \axi_wstrb_ns_i_i_a2_1[19]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_395, B => N_394, Y => N_523_1);
    
    \HADDR_sync[12]\ : SLE
      port map(D => HADDR_d(12), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12));
    
    \WDATA_i_i_o2[25]\ : CFG4
      generic map(INIT => x"6F0F")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \burstcount_reg[0]_net_1\, C => N_396, D => 
        \WDATA_i_i_o2_1[25]_net_1\, Y => N_390);
    
    \rdch_write_data_r[42]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(42), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[42]_net_1\);
    
    \un34_i_a2_0_a2_1[1]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \axi_wstrb[10]_net_1\, B => 
        \axi_wstrb[9]_net_1\, C => \axi_wstrb[6]_net_1\, Y => 
        \un34_i_a2_0_a2_1[1]_net_1\);
    
    \rdch_write_data_r[53]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(53), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[53]_net_1\);
    
    \burstcount_reg[3]\ : SLE
      port map(D => \SUM_i_m3[3]\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \burstcount_reg[3]_net_1\);
    
    \rdch_fifo_wr_data[30]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[62]_net_1\, B => 
        \rdch_write_data_r[30]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(30));
    
    \WDATA_i_o4_i_o2_RNIODKK3[4]\ : CFG4
      generic map(INIT => x"00D8")

      port map(A => N_396, B => N_435, C => N_428, D => 
        WDATA_sn_N_17_mux, Y => N_382_i);
    
    \WDATA_i_o2_i_RNISFMG3[31]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_223, B => N_215, C => WDATA_sn_N_17_mux, D
         => N_373, Y => N_202_i);
    
    \un34_i_a2_5_a2_1[4]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \axi_wstrb[19]_net_1\, B => 
        \axi_wstrb[18]_net_1\, C => \axi_wstrb[15]_net_1\, Y => 
        \un34_i_a2_5_a2_1[4]_net_1\);
    
    HWRITE_sync : SLE
      port map(D => HWRITE_d, CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \HWRITE_sync\);
    
    \HADDR_sync[26]\ : SLE
      port map(D => HADDR_d(26), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26));
    
    \axi_wstrb_ns_i_0_1[1]\ : CFG3
      generic map(INIT => x"DE")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_395, 
        Y => N_1723_1);
    
    \WDATA_1_m2_0_o2[58]\ : CFG4
      generic map(INIT => x"05CC")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \AWADDR_incr[2]_net_1\, C => N_397, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_140);
    
    \rdch_write_data_r[26]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(26), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[26]_net_1\);
    
    \HADDR_sync[24]\ : SLE
      port map(D => HADDR_d(24), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24));
    
    \un34_i_a2_5_a2_0[5]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \axi_wstrb[2]_net_1\, B => 
        \axi_wstrb[1]_net_1\, C => \axi_wstrb[0]_net_1\, Y => 
        N_550);
    
    \rdch_write_data_r[13]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(13), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[13]_net_1\);
    
    \axi_wstrb_ns_i_0_0[18]\ : CFG4
      generic map(INIT => x"4E5F")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => N_397, C => \axi_wstrb[7]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, Y => 
        \axi_wstrb_ns_i_0_0[18]_net_1\);
    
    \WDATA_i_i[26]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_414, B => N_417, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(26));
    
    wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_1_i_0_RNIOLJT : CFG4
      generic map(INIT => x"3331")

      port map(A => N_71_i_1, B => 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_1_i_0\, C => 
        \burstcount_reg[4]_net_1\, D => \burstcount_reg[3]_net_1\, 
        Y => N_71_i);
    
    \WDATA_i_i[25]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_413, B => N_416, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(25));
    
    \rdch_write_data_r[54]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(54), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[54]_net_1\);
    
    \rdch_write_data_r[25]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(25), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[25]_net_1\);
    
    \rdch_write_data_r[57]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(57), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[57]_net_1\);
    
    \rdch_write_data_r[30]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(30), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[30]_net_1\);
    
    \axi_current_state_ns_0[0]\ : CFG4
      generic map(INIT => x"FFCE")

      port map(A => \axi_current_state[0]_net_1\, B => 
        latch_wr_resp_set_xhdl66_0_sqmuxa, C => N_83, D => N_105, 
        Y => \axi_current_state_ns[0]\);
    
    \rdch_write_data_r[14]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(14), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[14]_net_1\);
    
    \rdch_fifo_wr_data[26]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[58]_net_1\, B => 
        \rdch_write_data_r[26]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(26));
    
    axi_read_data_xhdl68_1_i_i_a3 : CFG4
      generic map(INIT => x"8880")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_RVALID, B => 
        \axi_current_state[0]_net_1\, C => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_RREADY\, Y => 
        \axi_read_data_xhdl68_1_i_i_a3\);
    
    \AWADDR_incr_9_i_o2[2]\ : CFG4
      generic map(INIT => x"CCDF")

      port map(A => N_265, B => wready_m_xhdl2, C => 
        \AWADDR_incr[1]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_346);
    
    \rdch_fifo_wr_data[12]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[44]_net_1\, B => 
        \rdch_write_data_r[12]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(12));
    
    \WDATA_i_i[30]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_390, B => N_392, C => N_440, D => N_328, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(30));
    
    HADDR_sync_154 : CFG4
      generic map(INIT => x"E4F0")

      port map(A => \latch_ahb_sig_sync_d\, B => HADDR_d(1), C
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, D => 
        latch_ahb_sig_sync, Y => \HADDR_sync_154\);
    
    \rdch_fifo_wr_data[29]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[61]_net_1\, B => 
        \rdch_write_data_r[29]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(29));
    
    \rdch_write_data_r[17]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(17), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[17]_net_1\);
    
    \WDATA_i_i[18]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_420, B => N_424, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(18));
    
    \WDATA_1_0[49]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_423, B => N_140, C => N_139, D => N_419, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(49));
    
    \burstcount_reg[2]\ : SLE
      port map(D => N_69_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \burstcount_reg[2]_net_1\);
    
    \WDATA_0[33]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_194, B => N_159, C => N_150, D => N_142, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(33));
    
    \axi_current_state_ns_0_a3_1[0]\ : CFG4
      generic map(INIT => x"008A")

      port map(A => \axi_current_state[5]_net_1\, B => 
        ahb_rd_req_sync, C => \ahb_rd_req_sync_d\, D => 
        ahb_wr_done_sync, Y => N_105);
    
    \WDATA_0[43]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_291, B => N_194, C => N_142, D => N_284, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(43));
    
    \un34_i_a2_4_a2_2_RNI4P52[6]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \axi_wstrb[20]_net_1\, B => 
        \un34_i_a2_4_a2_2[6]_net_1\, C => \axi_wstrb[23]_net_1\, 
        D => \axi_wstrb[22]_net_1\, Y => N_1446_i);
    
    \WDATA_i_i[16]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_418, B => N_422, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(16));
    
    \HADDR_sync[8]\ : SLE
      port map(D => HADDR_d(8), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8));
    
    \rdch_write_data_r[2]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(2), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[2]_net_1\);
    
    \axi_wstrb_RNO[14]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[14]_net_1\, Y => 
        N_1727_i);
    
    \HADDR_sync[16]\ : SLE
      port map(D => HADDR_d(16), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16));
    
    ahb_rd_req_sync_d : SLE
      port map(D => ahb_rd_req_sync, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ahb_rd_req_sync_d\);
    
    \HADDR_sync[14]\ : SLE
      port map(D => HADDR_d(14), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14));
    
    \axi_wstrb[14]\ : SLE
      port map(D => N_1727_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[14]_net_1\);
    
    \WDATA_0_0[38]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_411, B => N_194, C => N_142, D => N_410, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(38));
    
    \rdch_write_data_r[32]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(32), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[32]_net_1\);
    
    \WDATA_i_o4_i_o2_RNIBTUD3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_281, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_288, Y => N_272_i);
    
    WRCH_fifo_rd_en_iv_i_o3 : CFG2
      generic map(INIT => x"7")

      port map(A => N_71_i, B => \burstcount_reg[0]_net_1\, Y => 
        N_98);
    
    \rdch_fifo_wr_data[15]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[47]_net_1\, B => 
        \rdch_write_data_r[15]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(15));
    
    \HSIZE_sync[1]\ : SLE
      port map(D => \HSIZE_sync_151\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\);
    
    wvalid_set_r_1_0_a3 : CFG2
      generic map(INIT => x"4")

      port map(A => \wvalid_reg\, B => \axi_current_state_2\, Y
         => wvalid_set_r_1);
    
    \un34_i_a2_4_a2_0[2]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \axi_wstrb[11]_net_1\, B => 
        \axi_wstrb[8]_net_1\, C => N_552, Y => N_563);
    
    \axi_wstrb[19]\ : SLE
      port map(D => N_1717_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[19]_net_1\);
    
    \axi_wstrb[18]\ : SLE
      port map(D => N_1719_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[18]_net_1\);
    
    \AWADDR_incr_9_i_m2[1]\ : CFG4
      generic map(INIT => x"AAC3")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, B
         => \AWADDR_incr[1]_net_1\, C => N_280, D => N_48_i, Y
         => \AWADDR_incr_9_i_m2[1]_net_1\);
    
    \axi_wstrb_RNO[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[2]_net_1\, Y => 
        N_1751_i);
    
    \burstcount_reg[1]\ : SLE
      port map(D => N_68_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \burstcount_reg[1]_net_1\);
    
    \axi_wstrb_RNO[16]\ : CFG4
      generic map(INIT => x"0D08")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \axi_wstrb[16]_net_1\, C => N_1723_1, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, Y => N_1723_i);
    
    \axi_wstrb_RNO[15]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[15]_net_1\, Y => 
        N_1725_i);
    
    \axi_wstrb[24]\ : SLE
      port map(D => N_1708_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[24]_net_1\);
    
    \axi_wstrb_ns_i_i[19]\ : CFG4
      generic map(INIT => x"C0EA")

      port map(A => N_551, B => \axi_wstrb[6]_net_1\, C => 
        N_523_1, D => N_397, Y => \axi_wstrb_ns_i_i[19]_net_1\);
    
    wvalid_reg_r_RNI3M6A1 : CFG4
      generic map(INIT => x"8000")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_WREADY, B => N_82, 
        C => \wvalid_reg_r\, D => \axi_current_state_2\, Y => 
        N_67_i_0);
    
    \rdch_write_data_r[60]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(60), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[60]_net_1\);
    
    \rdch_write_data_r[28]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(28), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[28]_net_1\);
    
    \axi_wstrb_ns_i_0_0[15]\ : CFG4
      generic map(INIT => x"33AF")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, B
         => \axi_wstrb[10]_net_1\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => 
        \axi_wstrb_ns_i_0_0[15]_net_1\);
    
    \WDATA_1_0[58]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_417, B => N_140, C => N_139, D => N_414, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(58));
    
    \un1_burstcount_reg_2_1.SUM_i_o3[3]\ : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \burstcount_reg[0]_net_1\, B => N_67_i_0, C
         => \burstcount_reg[2]_net_1\, D => 
        \burstcount_reg[1]_net_1\, Y => N_86);
    
    \WDATA_i_o4_i_o2_RNIQFKK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_286, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_293, Y => N_277_i);
    
    un1_axi_current_state_5_i_o3 : CFG2
      generic map(INIT => x"E")

      port map(A => \un1_axi_current_state_5_i_o3_sx\, B => 
        \burstcount_reg[0]_net_1\, Y => N_82);
    
    \axi_current_state_RNIPMOS1[3]\ : CFG4
      generic map(INIT => x"C8C0")

      port map(A => \burstcount_reg[0]_net_1\, B => 
        \axi_current_state_2\, C => \N_72_i\, D => N_71_i, Y => 
        N_73_i_0);
    
    \WDATA_1_0[56]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_425, B => N_140, C => N_139, D => N_421, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(56));
    
    \rdch_write_data_r[43]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(43), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[43]_net_1\);
    
    \axi_wstrb_ns_0_i_m2[3]\ : CFG4
      generic map(INIT => x"A8FD")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, D => N_395, Y
         => N_444);
    
    \rdch_write_data_r[21]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(21), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[21]_net_1\);
    
    \rdch_write_data_r[5]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(5), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[5]_net_1\);
    
    \HADDR_sync[7]\ : SLE
      port map(D => HADDR_d(7), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7));
    
    wvalid_reg_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => WLAST, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, Y => N_99_i);
    
    \rdch_fifo_wr_data[18]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[50]_net_1\, B => 
        \rdch_write_data_r[18]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(18));
    
    \rdch_write_data_r[7]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(7), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[7]_net_1\);
    
    \WDATA_i_o4_i_o2_RNINBJK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_148, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_157, Y => N_134_i);
    
    \WDATA_i_o2_i_RNINBNG3[31]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_221, B => N_213, C => WDATA_sn_N_17_mux, D
         => N_373, Y => N_200_i);
    
    \un34_i_a2_5_a2_2_RNIPV6O[3]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => \un34_i_a2_5_a2_2[3]_net_1\, B => N_563, C
         => \axi_wstrb[15]_net_1\, D => \axi_wstrb[14]_net_1\, Y
         => N_1449_i);
    
    rready_set_xhdl69_1_i_i_o3 : CFG2
      generic map(INIT => x"7")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_RVALID, B => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, Y => N_83);
    
    \WDATA_0[22]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_429, B => N_436, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(22));
    
    \axi_current_state[0]\ : SLE
      port map(D => \axi_current_state_ns[5]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state[0]_net_1\);
    
    \WDATA_0[35]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_194, B => N_157, C => N_148, D => N_142, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(35));
    
    \AWADDR_incr[2]\ : SLE
      port map(D => \AWADDR_incr_9_i_m2[2]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWADDR_incr[2]_net_1\);
    
    \WDATA_0[45]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_289, B => N_194, C => N_142, D => N_282, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(45));
    
    \axi_wstrb_RNO[0]\ : CFG4
      generic map(INIT => x"AA80")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \axi_wstrb[0]_net_1\, C => N_395, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_1755_i);
    
    \rdch_write_data_r[44]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(44), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[44]_net_1\);
    
    \rdch_fifo_wr_data[31]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[63]_net_1\, B => 
        \rdch_write_data_r[31]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(31));
    
    \WDATA_i_o2_i_m2[31]\ : CFG4
      generic map(INIT => x"5F88")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, D => 
        \WDATA_i_o2_i_m2_1[31]_net_1\, Y => N_330);
    
    \rdch_write_data_r[62]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(62), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[62]_net_1\);
    
    \axi_current_state[5]\ : SLE
      port map(D => \axi_current_state_ns[0]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state[5]_net_1\);
    
    \WDATA_i_i[24]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_421, B => N_425, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(24));
    
    \rdch_write_data_r[47]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(47), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[47]_net_1\);
    
    \WDATA_i_o2_i_RNISHOG3[31]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_218, B => N_210, C => WDATA_sn_N_17_mux, D
         => N_373, Y => N_197_i);
    
    \rdch_fifo_wr_data[10]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[42]_net_1\, B => 
        \rdch_write_data_r[10]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(10));
    
    \gen_start_for_rdch_read.axi_read_rlast_xhdl26_1_0_a3\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_83, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_RREADY\, Y => 
        axi_read_rlast_xhdl26_1);
    
    \WDATA_i_o4_i_o2_RNIL9JK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_149, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_158, Y => N_135_i);
    
    \un34_i_a2_5_a2_1_RNIRV3N[4]\ : CFG4
      generic map(INIT => x"FFF7")

      port map(A => \un34_i_a2_5_a2_1[4]_net_1\, B => N_563, C
         => \axi_wstrb[17]_net_1\, D => \axi_wstrb[14]_net_1\, Y
         => N_1448_i);
    
    \HADDR_sync[25]\ : SLE
      port map(D => HADDR_d(25), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25));
    
    \axi_wstrb_RNO[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[1]_net_1\, Y => 
        N_1753_i);
    
    awaddr_awvalid_clr_d_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \axi_current_state_3\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, Y => N_88_i);
    
    \WDATA_i_o4_i_o2_RNIRFJK3[4]\ : CFG4
      generic map(INIT => x"00D8")

      port map(A => N_396, B => N_433, C => N_426, D => 
        WDATA_sn_N_17_mux, Y => N_380_i);
    
    \axi_wstrb_ns_i_0_o2[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, Y => N_395);
    
    axi_read_rlast_xhdl26 : SLE
      port map(D => axi_read_rlast_xhdl26_1, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        axi_read_rlast);
    
    \rdch_write_data_r[56]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(56), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[56]_net_1\);
    
    store_ahb_sig : CFG2
      generic map(INIT => x"2")

      port map(A => latch_ahb_sig_sync, B => 
        \latch_ahb_sig_sync_d\, Y => \store_ahb_sig\);
    
    HSIZE_sync_151 : CFG4
      generic map(INIT => x"E4F0")

      port map(A => \latch_ahb_sig_sync_d\, B => HSIZE_d(1), C
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, D => 
        latch_ahb_sig_sync, Y => \HSIZE_sync_151\);
    
    \un34_i_a2_4_a2_2[6]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \axi_wstrb[17]_net_1\, B => 
        \axi_wstrb[1]_net_1\, C => \axi_wstrb[0]_net_1\, D => 
        \axi_wstrb[14]_net_1\, Y => \un34_i_a2_4_a2_2[6]_net_1\);
    
    \axi_wstrb_ns_i_0_m2[2]\ : CFG4
      generic map(INIT => x"F011")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, C => 
        \axi_wstrb[23]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, Y => N_443);
    
    wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_i_0_RNICFBE : CFG2
      generic map(INIT => x"2")

      port map(A => N_82, B => 
        \wrch_fifo_rd_en_xhdl22_xhdl65_1_sqmuxa_i_0\, Y => 
        \N_72_i\);
    
    \WDATA_1[53]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_221, B => N_140, C => N_139, D => N_213, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(53));
    
    \rdch_fifo_wr_data[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[32]_net_1\, B => 
        \rdch_write_data_r[0]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(0));
    
    \un1_burstcount_reg_2_1.N_69_i\ : CFG3
      generic map(INIT => x"09")

      port map(A => N_91, B => \burstcount_reg[2]_net_1\, C => 
        N_79, Y => N_69_i);
    
    \rdch_write_data_r[55]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(55), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[55]_net_1\);
    
    \rdch_write_data_r[16]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(16), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[16]_net_1\);
    
    \WDATA_0[41]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_293, B => N_194, C => N_142, D => N_286, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(41));
    
    HMASTLOCK_sync : SLE
      port map(D => HMASTLOCK_d, CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0);
    
    \HADDR_sync[19]\ : SLE
      port map(D => HADDR_d(19), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19));
    
    \rdch_write_data_r[33]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(33), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[33]_net_1\);
    
    \un34_i_a2_5_a2_2[3]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \axi_wstrb[16]_net_1\, B => 
        \axi_wstrb[12]_net_1\, C => \axi_wstrb[4]_net_1\, Y => 
        \un34_i_a2_5_a2_2[3]_net_1\);
    
    \WDATA_i_o4_i_o2_RNIPDJK3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_147, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_156, Y => N_133_i);
    
    \axi_current_state[4]\ : SLE
      port map(D => \axi_current_state_ns[1]\, CLK => SDRCLK_c, 
        EN => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \axi_current_state_3\);
    
    \WDATA_1_o2_0_o2_0[58]\ : CFG3
      generic map(INIT => x"25")

      port map(A => \burstcount_reg[0]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, Y => N_389);
    
    rready_set_xhdl69_1_i_i : CFG3
      generic map(INIT => x"EA")

      port map(A => \axi_current_state_0\, B => N_83, C => 
        \axi_current_state[0]_net_1\, Y => 
        \rready_set_xhdl69_1_i_i\);
    
    \rdch_write_data_r[4]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(4), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[4]_net_1\);
    
    \rdch_fifo_wr_data[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[35]_net_1\, B => 
        \rdch_write_data_r[3]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(3));
    
    \swap_rd_data_byte[2]\ : SLE
      port map(D => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, CLK
         => SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \swap_rd_data_byte[2]_net_1\);
    
    \rdch_fifo_wr_data[22]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[54]_net_1\, B => 
        \rdch_write_data_r[22]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(22));
    
    un1_axi_current_state_5_i_o3_sx : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \burstcount_reg[4]_net_1\, B => 
        \burstcount_reg[3]_net_1\, C => \burstcount_reg[2]_net_1\, 
        D => \burstcount_reg[1]_net_1\, Y => 
        \un1_axi_current_state_5_i_o3_sx\);
    
    \rdch_write_data_r[29]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(29), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[29]_net_1\);
    
    \rdch_write_data_r[15]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(15), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[15]_net_1\);
    
    \WDATA_i_o4_i_o2_RNITHJK3[4]\ : CFG4
      generic map(INIT => x"00D8")

      port map(A => N_396, B => N_411, C => N_410, D => 
        WDATA_sn_N_17_mux, Y => N_278_i);
    
    \araddr_arvalid_clr_d\ : SLE
      port map(D => N_274_i_0, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        araddr_arvalid_clr_d_net_1);
    
    WLAST_0_a2_RNO : CFG4
      generic map(INIT => x"FFBF")

      port map(A => \axi_current_state_0\, B => \wvalid_reg\, C
         => \wvalid_reg_r\, D => \axi_current_state[0]_net_1\, Y
         => N_100_i);
    
    WLAST_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => N_100_i, B => un1_axi_current_state_i, Y => 
        WLAST);
    
    \axi_wstrb_RNO[24]\ : CFG4
      generic map(INIT => x"080D")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, B
         => \axi_wstrb[24]_net_1\, C => N_1723_1, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, Y => N_1708_i);
    
    \axi_wstrb_ns_i_0_m2[13]\ : CFG4
      generic map(INIT => x"BB0F")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, C => 
        \axi_wstrb[12]_net_1\, D => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => N_446);
    
    \rdch_write_data_r[34]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(34), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[34]_net_1\);
    
    \WDATA_1_0[48]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_422, B => N_140, C => N_139, D => N_418, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(48));
    
    HSIZE_sync_150 : CFG4
      generic map(INIT => x"E4F0")

      port map(A => \latch_ahb_sig_sync_d\, B => HSIZE_d(0), C
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, D => 
        latch_ahb_sig_sync, Y => \HSIZE_sync_150\);
    
    \axi_wstrb[1]\ : SLE
      port map(D => N_1753_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[1]_net_1\);
    
    \HADDR_sync[15]\ : SLE
      port map(D => HADDR_d(15), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15));
    
    \rdch_write_data_r[37]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(37), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[37]_net_1\);
    
    \HADDR_sync[6]\ : SLE
      port map(D => HADDR_d(6), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6));
    
    \axi_wstrb_RNO[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[11]_net_1\, Y => 
        N_1733_i);
    
    \rdch_fifo_wr_data[17]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[49]_net_1\, B => 
        \rdch_write_data_r[17]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(17));
    
    \axi_wstrb[16]\ : SLE
      port map(D => N_1723_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[16]_net_1\);
    
    \awaddr_awvalid_clr_d\ : SLE
      port map(D => N_88_i, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        awaddr_awvalid_clr_d_net_1);
    
    \rdch_fifo_wr_data[25]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[57]_net_1\, B => 
        \rdch_write_data_r[25]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(25));
    
    \WDATA_i_o4_i_o2_RNI9RUD3[4]\ : CFG4
      generic map(INIT => x"2320")

      port map(A => N_282, B => WDATA_sn_N_17_mux, C => N_396, D
         => N_289, Y => N_273_i);
    
    \rdch_fifo_wr_data[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[33]_net_1\, B => 
        \rdch_write_data_r[1]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(1));
    
    \WDATA_0[32]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_194, B => N_160, C => N_151, D => N_142, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(32));
    
    \AWADDR_incr_9_i_o2[1]\ : CFG4
      generic map(INIT => x"F7FF")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_WVALID\, B => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, D => N_265, Y
         => N_280);
    
    \WDATA_0[27]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => N_431, B => N_438, C => N_392, D => N_390, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(27));
    
    \WDATA_0[42]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_292, B => N_194, C => N_142, D => N_285, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(42));
    
    \AWADDR_incr[0]\ : SLE
      port map(D => \AWADDR_incr_9_i_m2[0]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWADDR_incr[0]_net_1\);
    
    \WDATA_i_o2_i_RNIL9NG3[31]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_222, B => N_214, C => WDATA_sn_N_17_mux, D
         => N_373, Y => N_201_i);
    
    \rdch_write_data_r[63]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(63), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[63]_net_1\);
    
    \WDATA_1[55]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_437, B => N_140, C => N_139, D => N_430, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(55));
    
    \rdch_write_data_r[58]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(58), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[58]_net_1\);
    
    \rdch_write_data_r[0]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(0), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[0]_net_1\);
    
    \un34_i_a2_5_a2_2[5]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \axi_wstrb[21]_net_1\, B => 
        \axi_wstrb[20]_net_1\, C => \axi_wstrb[18]_net_1\, D => 
        \axi_wstrb[11]_net_1\, Y => \un34_i_a2_5_a2_2[5]_net_1\);
    
    un43_hburst_sync_i_i : CFG3
      generic map(INIT => x"20")

      port map(A => \axi_current_state_3\, B => 
        awaddr_awvalid_clr_d_net_1, C => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, Y => N_48_i);
    
    \WDATA_1[63]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_217, B => N_140, C => N_139, D => N_209, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(63));
    
    \rdch_fifo_wr_data[13]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[45]_net_1\, B => 
        \rdch_write_data_r[13]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(13));
    
    wvalid_clr_t : SLE
      port map(D => WLAST, CLK => SDRCLK_c, EN => VCC_net_1, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \wvalid_clr_t\);
    
    \WDATA_0[36]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_194, B => N_156, C => N_147, D => N_142, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(36));
    
    \rdch_write_data_r[51]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(51), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[51]_net_1\);
    
    \rdch_write_data_r[18]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(18), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[18]_net_1\);
    
    \AWADDR_incr_9_i_o2_0[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \AWADDR_incr[0]_net_1\, Y => N_265);
    
    \WDATA_0[46]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_288, B => N_194, C => N_142, D => N_281, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(46));
    
    \rdch_fifo_wr_data[28]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[60]_net_1\, B => 
        \rdch_write_data_r[28]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(28));
    
    \rdch_write_data_r[46]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(46), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[46]_net_1\);
    
    \rdch_write_data_r[11]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(11), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[11]_net_1\);
    
    \rdch_write_data_r[9]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(9), CLK => 
        SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn => 
        ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[9]_net_1\);
    
    \rdch_fifo_wr_data[11]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[43]_net_1\, B => 
        \rdch_write_data_r[11]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(11));
    
    \axi_wstrb_RNO[19]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \axi_wstrb_ns_i_0_0[6]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, C => N_395, Y
         => N_1717_i);
    
    \WDATA_i_o2_i_m2_1[31]\ : CFG3
      generic map(INIT => x"35")

      port map(A => \AWADDR_incr[2]_net_1\, B => 
        \burstcount_reg[0]_net_1\, C => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, Y => 
        \WDATA_i_o2_i_m2_1[31]_net_1\);
    
    HADDR_sync_153 : CFG4
      generic map(INIT => x"E2F0")

      port map(A => HADDR_d(0), B => \latch_ahb_sig_sync_d\, C
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, D => 
        latch_ahb_sig_sync, Y => \HADDR_sync_153\);
    
    \un34_i_a2_0_a2_1[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \axi_wstrb[4]_net_1\, B => 
        \axi_wstrb[5]_net_1\, Y => N_558);
    
    \rdch_write_data_r[45]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(45), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[45]_net_1\);
    
    \AWADDR_incr[1]\ : SLE
      port map(D => \AWADDR_incr_9_i_m2[1]_net_1\, CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \AWADDR_incr[1]_net_1\);
    
    \axi_wstrb_RNO[4]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \axi_wstrb[4]_net_1\, B => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, C => N_394, D
         => N_395, Y => N_1747_i);
    
    \axi_wstrb_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_523_1, B => \axi_wstrb[5]_net_1\, Y => 
        N_1745_i);
    
    \un1_burstcount_reg_2_1.N_68_i\ : CFG4
      generic map(INIT => x"5014")

      port map(A => N_79, B => N_67_i_0, C => 
        \burstcount_reg[1]_net_1\, D => \burstcount_reg[0]_net_1\, 
        Y => N_68_i);
    
    \WDATA_1[51]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_223, B => N_140, C => N_139, D => N_215, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(51));
    
    \rdch_fifo_wr_data[20]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[52]_net_1\, B => 
        \rdch_write_data_r[20]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(20));
    
    un1_rd_data_c_xhdl44_1_sqmuxa_i : CFG4
      generic map(INIT => x"F0F4")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, C => 
        \un1_rd_data_c_xhdl44_1_sqmuxa_i_0\, D => N_395, Y => 
        N_384);
    
    \WDATA_1_o2_0_o2[58]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => N_389, C => N_194, Y => N_139);
    
    \axi_wstrb_RNO[10]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, B
         => \axi_wstrb_ns_i_0_0[15]_net_1\, C => N_395, Y => 
        N_1735_i);
    
    \WDATA_0[40]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_435, B => N_194, C => N_142, D => N_428, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(40));
    
    \rdch_write_data_r[20]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(20), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[20]_net_1\);
    
    \rdch_fifo_wr_data[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[36]_net_1\, B => 
        \rdch_write_data_r[4]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(4));
    
    \HADDR_sync[21]\ : SLE
      port map(D => HADDR_d(21), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21));
    
    \un34_i_a2_4_a2_0_0[2]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \axi_wstrb[9]_net_1\, B => 
        \axi_wstrb[13]_net_1\, Y => \un34_i_a2_4_a2_0[2]_net_1\);
    
    \axi_current_state_ns_0_o3[5]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => COREAHBLTOAXI_0_AXIMasterIF_AWREADY, B => 
        \axi_current_state_3\, C => N_274_i_0, Y => N_81);
    
    \HADDR_sync[5]\ : SLE
      port map(D => HADDR_d(5), CLK => SDRCLK_c, EN => 
        \store_ahb_sig\, ALn => ARESET_n, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5));
    
    \WDATA_1_0[50]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_424, B => N_140, C => N_139, D => N_420, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(50));
    
    latch_ahb_sig_sync_d : SLE
      port map(D => latch_ahb_sig_sync, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \latch_ahb_sig_sync_d\);
    
    \axi_wstrb[7]\ : SLE
      port map(D => N_1741_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[7]_net_1\);
    
    \HADDR_sync[2]\ : SLE
      port map(D => \HADDR_sync_155\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\);
    
    wvalid_reg : SLE
      port map(D => N_99_i, CLK => SDRCLK_c, EN => 
        \wvalid_reg_1_sqmuxa_i_0\, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wvalid_reg\);
    
    un1_rd_data_c_xhdl44_1_sqmuxa_i_x2 : CFG2
      generic map(INIT => x"6")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[0]\, Y => N_555);
    
    \axi_wstrb[13]\ : SLE
      port map(D => N_1729_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[13]_net_1\);
    
    \HSIZE_sync[0]\ : SLE
      port map(D => \HSIZE_sync_150\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\);
    
    \rdch_fifo_wr_data[14]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[46]_net_1\, B => 
        \rdch_write_data_r[14]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(14));
    
    \axi_wstrb[17]\ : SLE
      port map(D => N_1721_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[17]_net_1\);
    
    \rdch_fifo_wr_data[9]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[41]_net_1\, B => 
        \rdch_write_data_r[9]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(9));
    
    \axi_wstrb_ns_i_0_o2[18]\ : CFG2
      generic map(INIT => x"7")

      port map(A => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, B
         => \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, Y => N_397);
    
    \axi_current_state_ns_o2_0_o3[2]\ : CFG4
      generic map(INIT => x"EAC0")

      port map(A => \axi_current_state_2\, B => \HWRITE_sync\, C
         => N_81, D => N_82, Y => \axi_current_state_ns[2]\);
    
    \rdch_write_data_r[36]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(36), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[36]_net_1\);
    
    \rdch_write_data_r[59]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(59), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[59]_net_1\);
    
    \rdch_write_data_r[48]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(48), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[48]_net_1\);
    
    \WDATA_0[37]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_433, B => N_194, C => N_142, D => N_426, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(37));
    
    \axi_wstrb[23]\ : SLE
      port map(D => N_1710_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[23]_net_1\);
    
    \axi_wstrb[0]\ : SLE
      port map(D => N_1755_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[0]_net_1\);
    
    \rdch_write_data_r[22]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(22), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[22]_net_1\);
    
    awaddr_awvalid_clr_d_RNIL7OF : CFG2
      generic map(INIT => x"2")

      port map(A => \axi_current_state_3\, B => 
        awaddr_awvalid_clr_d_net_1, Y => N_75_i);
    
    \WDATA_1[52]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => N_222, B => N_140, C => N_139, D => N_214, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(52));
    
    \axi_wstrb[5]\ : SLE
      port map(D => N_1745_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \axi_wstrb[5]_net_1\);
    
    \rdch_fifo_wr_data[5]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \rdch_write_data_r[37]_net_1\, B => 
        \rdch_write_data_r[5]_net_1\, C => N_384, Y => 
        rdch_fifo_wr_data(5));
    
    \rdch_write_data_r[35]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(35), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[35]_net_1\);
    
    \un34_i_a2_0_a2_1_RNIAE571[1]\ : CFG4
      generic map(INIT => x"F7FF")

      port map(A => \un34_i_a2_0_a2_1[1]_net_1\, B => N_552, C
         => \axi_wstrb[8]_net_1\, D => N_558, Y => N_1451_i);
    
    \rdch_write_data_r[41]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(41), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[41]_net_1\);
    
    \rdch_write_data_r[19]\ : SLE
      port map(D => COREAHBLTOAXI_0_AXIMasterIF_RDATA(19), CLK
         => SDRCLK_c, EN => \axi_read_data_xhdl68_1_i_i_a3\, ALn
         => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rdch_write_data_r[19]_net_1\);
    
    \axi_wstrb_RNIC8H11[7]\ : CFG4
      generic map(INIT => x"EFFF")

      port map(A => \axi_wstrb[7]_net_1\, B => 
        \axi_wstrb[6]_net_1\, C => N_558, D => N_552, Y => 
        N_1452_i);
    
    \WDATA_0[34]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_194, B => N_158, C => N_149, D => N_142, Y
         => COREAHBLTOAXI_0_AXIMasterIF_WDATA(34));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAHBLtoAXI_AHBAccessControlHX is

    port( CoreAHBLite_0_AHBmslave10_HADDR     : in    std_logic_vector(27 downto 0);
          HADDR_d                             : out   std_logic_vector(27 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE     : in    std_logic_vector(1 downto 0);
          HSIZE_d                             : out   std_logic_vector(1 downto 0);
          rdch_read_data                      : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HRDATA    : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA    : in    std_logic_vector(31 downto 0);
          wrch_hwdata_r                       : out   std_logic_vector(31 downto 0);
          xhdl1222_0                          : in    std_logic;
          synchronizer_1_0                    : in    std_logic;
          masterAddrInProg_0                  : in    std_logic;
          current_state_0                     : out   std_logic;
          N_92                                : in    std_logic;
          m0PrevDataSlaveReady                : in    std_logic;
          N_91                                : in    std_logic;
          post_sync_1_reg                     : in    std_logic;
          rdch_fifo_empty                     : in    std_logic;
          N_163_i                             : out   std_logic;
          hsel2                               : in    std_logic;
          hsel2_0_a2_1                        : in    std_logic;
          valid_ahbcmd_i_o3_1                 : out   std_logic;
          rdch_fifo_rd_en_r                   : out   std_logic;
          latch_ahb_sig                       : out   std_logic;
          BVALID_sync                         : in    std_logic;
          ahb_wr_done                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK : in    std_logic;
          HMASTLOCK_d                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE    : in    std_logic;
          HWRITE_d                            : out   std_logic;
          SDRCLK_c                            : in    std_logic;
          ARESET_n                            : in    std_logic;
          ahb_busyidle_cyc_i                  : out   std_logic;
          ahb_busyidle_cyc                    : out   std_logic
        );

end CoreAHBLtoAXI_AHBAccessControlHX;

architecture DEF_ARCH of CoreAHBLtoAXI_AHBAccessControlHX is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \ahb_busyidle_cyc\, \HTRANS_d_xhdl16[1]_net_1\, 
        \HTRANS_d_xhdl16_i[1]\, VCC_net_1, GND_net_1, 
        \wait_count_xhdl31[0]_net_1\, \wait_count_xhdl31_2[0]\, 
        \wait_count_xhdl31[1]_net_1\, N_141_i, 
        \rdch_fifo_rd_en_r_d\, latchahbcmd_xhdl34_1, 
        \current_state[1]_net_1\, \current_state[4]_net_1\, 
        \current_state[0]_net_1\, \current_state_ns[7]\, 
        \current_state_0\, N_149_i, \ahb_wr_done\, N_151_i, 
        \current_state[5]_net_1\, \current_state_ns[2]\, 
        \current_state_ns[3]\, \current_state[2]_net_1\, 
        \current_state_ns[5]\, \BVALID_sync_d\, 
        \rdch_fifo_rd_en_r\, N_335_i, 
        \current_state_ns_i_0_o2[1]_net_1\, burst_m2_0_a2_1, 
        burst_m2_0_a2_2, N_149_i_1, valid_ahbcmd_i_o3_1_net_1, 
        un1_current_state_2_i, fifo_rd_en_xhdl40_1_sqmuxa, N_357, 
        N_359, current_m2_e_0_1 : std_logic;

begin 

    current_state_0 <= \current_state_0\;
    valid_ahbcmd_i_o3_1 <= valid_ahbcmd_i_o3_1_net_1;
    rdch_fifo_rd_en_r <= \rdch_fifo_rd_en_r\;
    ahb_wr_done <= \ahb_wr_done\;
    ahb_busyidle_cyc <= \ahb_busyidle_cyc\;

    \hwdata_r_xhdl4[7]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(7), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(7));
    
    \HADDR_d_xhdl13[15]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(15), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(15));
    
    \RD_DATA_d1[10]\ : SLE
      port map(D => rdch_read_data(10), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(10));
    
    rdch_fifo_rd_en_r_xhdl6 : SLE
      port map(D => N_335_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rdch_fifo_rd_en_r\);
    
    \hwdata_r_xhdl4[4]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(4), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(4));
    
    latch_ahb_sig_xhdl9 : SLE
      port map(D => latchahbcmd_xhdl34_1, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        latch_ahb_sig);
    
    \HSIZE_d_xhdl17[0]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HSIZE(0), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HSIZE_d(0));
    
    BVALID_sync_d : SLE
      port map(D => BVALID_sync, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \BVALID_sync_d\);
    
    HMASTLOCK_d_xhdl19 : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HMASTLOCK, CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HMASTLOCK_d);
    
    \hwdata_r_xhdl4[10]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(10), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(10));
    
    \RD_DATA_d1[22]\ : SLE
      port map(D => rdch_read_data(22), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(22));
    
    \hwdata_r_xhdl4[17]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(17), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(17));
    
    un1_current_state_2_0_o2_RNIBD6G : CFG3
      generic map(INIT => x"01")

      port map(A => un1_current_state_2_i, B => 
        \current_state[2]_net_1\, C => \ahb_wr_done\, Y => 
        burst_m2_0_a2_1);
    
    \RD_DATA_d1[12]\ : SLE
      port map(D => rdch_read_data(12), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(12));
    
    \current_state_ns_0[5]\ : CFG4
      generic map(INIT => x"AEAA")

      port map(A => N_359, B => current_m2_e_0_1, C => 
        valid_ahbcmd_i_o3_1_net_1, D => masterAddrInProg_0, Y => 
        \current_state_ns[5]\);
    
    \RD_DATA_d1[21]\ : SLE
      port map(D => rdch_read_data(21), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(21));
    
    \HADDR_d_xhdl13[6]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(6), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(6));
    
    \HADDR_d_xhdl13[7]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(7), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(7));
    
    \RD_DATA_d1[4]\ : SLE
      port map(D => rdch_read_data(4), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(4));
    
    \hwdata_r_xhdl4[13]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(13), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(13));
    
    \valid_ahbcmd_i_o3_1\ : CFG4
      generic map(INIT => x"37FF")

      port map(A => m0PrevDataSlaveReady, B => N_92, C => 
        xhdl1222_0, D => \current_state_0\, Y => 
        valid_ahbcmd_i_o3_1_net_1);
    
    \RD_DATA_d1[11]\ : SLE
      port map(D => rdch_read_data(11), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(11));
    
    \hwdata_r_xhdl4[29]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(29), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(29));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \hwdata_r_xhdl4[1]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(1), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(1));
    
    \hwdata_r_xhdl4[16]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(16), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(16));
    
    HWRITE_d_xhdl14 : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWRITE, CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HWRITE_d);
    
    \hwdata_r_xhdl4[31]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(31), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(31));
    
    \HADDR_d_xhdl13[8]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(8), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(8));
    
    \HADDR_d_xhdl13[24]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(24), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(24));
    
    \HADDR_d_xhdl13[2]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(2), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(2));
    
    \current_state[1]\ : SLE
      port map(D => \current_state[4]_net_1\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \current_state[1]_net_1\);
    
    \HADDR_d_xhdl13[14]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(14), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(14));
    
    \RD_DATA_d1[24]\ : SLE
      port map(D => rdch_read_data(24), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(24));
    
    \current_state[2]\ : SLE
      port map(D => \current_state_ns[5]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \current_state[2]_net_1\);
    
    \wait_count_xhdl31_RNO[1]\ : CFG3
      generic map(INIT => x"48")

      port map(A => \wait_count_xhdl31[1]_net_1\, B => 
        \current_state[0]_net_1\, C => 
        \wait_count_xhdl31[0]_net_1\, Y => N_141_i);
    
    \RD_DATA_d1[23]\ : SLE
      port map(D => rdch_read_data(23), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(23));
    
    \hwdata_r_xhdl4[8]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(8), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(8));
    
    \HADDR_d_xhdl13[22]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(22), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(22));
    
    \HADDR_d_xhdl13[27]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(27), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(27));
    
    \hwdata_r_xhdl4[20]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(20), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(20));
    
    \hwdata_r_xhdl4[12]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(12), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(12));
    
    \HADDR_d_xhdl13[12]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(12), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(12));
    
    \current_state_ns_i_0_o2[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => \BVALID_sync_d\, B => \current_state_0\, C
         => \current_state[5]_net_1\, Y => 
        \current_state_ns_i_0_o2[1]_net_1\);
    
    \wait_count_xhdl31[0]\ : SLE
      port map(D => \wait_count_xhdl31_2[0]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wait_count_xhdl31[0]_net_1\);
    
    \RD_DATA_d1[14]\ : SLE
      port map(D => rdch_read_data(14), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(14));
    
    \hwdata_r_xhdl4[27]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(27), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(27));
    
    \HADDR_d_xhdl13[17]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(17), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(17));
    
    un1_current_state_2_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \current_state[4]_net_1\, B => 
        \current_state[0]_net_1\, Y => un1_current_state_2_i);
    
    \RD_DATA_d1[8]\ : SLE
      port map(D => rdch_read_data(8), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(8));
    
    \RD_DATA_d1[13]\ : SLE
      port map(D => rdch_read_data(13), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(13));
    
    \HTRANS_d_xhdl16[1]\ : SLE
      port map(D => VCC_net_1, CLK => SDRCLK_c, EN => 
        latchahbcmd_xhdl34_1, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \HTRANS_d_xhdl16[1]_net_1\);
    
    ahb_busyidle_cyc_xhdl21_RNIOAG6 : CFG1
      generic map(INIT => "01")

      port map(A => \ahb_busyidle_cyc\, Y => ahb_busyidle_cyc_i);
    
    \RD_DATA_d1[1]\ : SLE
      port map(D => rdch_read_data(1), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(1));
    
    \hwdata_r_xhdl4[14]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(14), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(14));
    
    \hwdata_r_xhdl4[5]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(5), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(5));
    
    \current_state[4]\ : SLE
      port map(D => \current_state_ns[3]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \current_state[4]_net_1\);
    
    \RD_DATA_d1[30]\ : SLE
      port map(D => rdch_read_data(30), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(30));
    
    \RD_DATA_d1[0]\ : SLE
      port map(D => rdch_read_data(0), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(0));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \wait_count_xhdl31[1]\ : SLE
      port map(D => N_141_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wait_count_xhdl31[1]_net_1\);
    
    \hwdata_r_xhdl4[15]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(15), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(15));
    
    \hwdata_r_xhdl4[23]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(23), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(23));
    
    \current_state[0]\ : SLE
      port map(D => \current_state_ns[7]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \current_state[0]_net_1\);
    
    \wait_count_xhdl31_2_a3_0_a2[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \current_state[0]_net_1\, B => 
        \wait_count_xhdl31[0]_net_1\, Y => 
        \wait_count_xhdl31_2[0]\);
    
    \current_state_RNI6Q721[5]\ : CFG3
      generic map(INIT => x"A2")

      port map(A => burst_m2_0_a2_1, B => 
        \current_state[5]_net_1\, C => \BVALID_sync_d\, Y => 
        burst_m2_0_a2_2);
    
    \hwdata_r_xhdl4[26]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(26), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(26));
    
    \HADDR_d_xhdl13[5]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(5), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(5));
    
    \RD_DATA_d1[27]\ : SLE
      port map(D => rdch_read_data(27), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(27));
    
    \hwdata_r_xhdl4[18]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(18), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(18));
    
    \HADDR_d_xhdl13[4]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(4), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(4));
    
    \HADDR_d_xhdl13[1]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(1), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(1));
    
    \RD_DATA_d1[26]\ : SLE
      port map(D => rdch_read_data(26), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(26));
    
    \RD_DATA_d1[25]\ : SLE
      port map(D => rdch_read_data(25), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(25));
    
    \RD_DATA_d1[17]\ : SLE
      port map(D => rdch_read_data(17), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(17));
    
    \hwdata_r_xhdl4[22]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(22), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(22));
    
    \RD_DATA_d1[16]\ : SLE
      port map(D => rdch_read_data(16), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(16));
    
    \RD_DATA_d1[15]\ : SLE
      port map(D => rdch_read_data(15), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(15));
    
    \HADDR_d_xhdl13[23]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(23), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(23));
    
    valid_ahbcmd_i_o3_1_RNITATE4 : CFG3
      generic map(INIT => x"02")

      port map(A => hsel2, B => valid_ahbcmd_i_o3_1_net_1, C => 
        CoreAHBLite_0_AHBmslave10_HWRITE, Y => N_163_i);
    
    \hwdata_r_xhdl4[0]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(0), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(0));
    
    \RD_DATA_d1[31]\ : SLE
      port map(D => rdch_read_data(31), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(31));
    
    \hwdata_r_xhdl4[24]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(24), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(24));
    
    \HADDR_d_xhdl13[13]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(13), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(13));
    
    \hwdata_r_xhdl4[6]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(6), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(6));
    
    \current_state_RNO_0[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => valid_ahbcmd_i_o3_1_net_1, B => hsel2_0_a2_1, 
        Y => N_149_i_1);
    
    \current_state[5]\ : SLE
      port map(D => \current_state_ns[2]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \current_state[5]_net_1\);
    
    \RD_DATA_d1[9]\ : SLE
      port map(D => rdch_read_data(9), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(9));
    
    \RD_DATA_d1[29]\ : SLE
      port map(D => rdch_read_data(29), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(29));
    
    \hwdata_r_xhdl4[11]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(11), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(11));
    
    valid_ahbcmd_i_o3_1_RNIQLPS4 : CFG4
      generic map(INIT => x"0080")

      port map(A => burst_m2_0_a2_2, B => hsel2_0_a2_1, C => 
        masterAddrInProg_0, D => valid_ahbcmd_i_o3_1_net_1, Y => 
        latchahbcmd_xhdl34_1);
    
    \hwdata_r_xhdl4[30]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(30), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(30));
    
    \hwdata_r_xhdl4[2]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(2), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(2));
    
    \HADDR_d_xhdl13[20]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(20), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(20));
    
    \current_state[6]\ : SLE
      port map(D => N_151_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \ahb_wr_done\);
    
    \RD_DATA_d1[2]\ : SLE
      port map(D => rdch_read_data(2), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(2));
    
    \hwdata_r_xhdl4[3]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(3), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(3));
    
    fifo_rd_en_xhdl40_1_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"02")

      port map(A => \wait_count_xhdl31_2[0]\, B => 
        rdch_fifo_empty, C => \wait_count_xhdl31[1]_net_1\, Y => 
        fifo_rd_en_xhdl40_1_sqmuxa);
    
    \RD_DATA_d1[19]\ : SLE
      port map(D => rdch_read_data(19), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(19));
    
    \HADDR_d_xhdl13[10]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(10), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(10));
    
    \current_state_ns_0[2]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => \BVALID_sync_d\, B => \ahb_wr_done\, C => 
        \current_state[5]_net_1\, Y => \current_state_ns[2]\);
    
    \hwdata_r_xhdl4[25]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(25), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(25));
    
    \HADDR_d_xhdl13[26]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(26), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(26));
    
    \RD_DATA_d1[5]\ : SLE
      port map(D => rdch_read_data(5), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(5));
    
    \HADDR_d_xhdl13[21]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(21), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(21));
    
    \current_state_ns_0_RNO[5]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \current_state_ns_i_0_o2[1]_net_1\, B => 
        hsel2_0_a2_1, C => N_91, Y => current_m2_e_0_1);
    
    \HADDR_d_xhdl13[9]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(9), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(9));
    
    \HADDR_d_xhdl13[16]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(16), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(16));
    
    \RD_DATA_d1[6]\ : SLE
      port map(D => rdch_read_data(6), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(6));
    
    \HADDR_d_xhdl13[11]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(11), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(11));
    
    \HADDR_d_xhdl13[3]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(3), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(3));
    
    \RD_DATA_d1[3]\ : SLE
      port map(D => rdch_read_data(3), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(3));
    
    ahb_busyidle_cyc_xhdl21 : SLE
      port map(D => \HTRANS_d_xhdl16_i[1]\, CLK => SDRCLK_c, EN
         => VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ahb_busyidle_cyc\);
    
    \current_state_RNO[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAHBLite_0_AHBmslave10_HWRITE, B => 
        valid_ahbcmd_i_o3_1_net_1, Y => N_151_i);
    
    \current_state_ns_0_a2_0[7]\ : CFG3
      generic map(INIT => x"28")

      port map(A => \current_state[2]_net_1\, B => 
        synchronizer_1_0, C => post_sync_1_reg, Y => N_357);
    
    \current_state[7]\ : SLE
      port map(D => N_149_i, CLK => SDRCLK_c, EN => VCC_net_1, 
        ALn => ARESET_n, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \current_state_0\);
    
    \hwdata_r_xhdl4[28]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(28), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(28));
    
    \current_state_ns_a3_0_a2[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \wait_count_xhdl31_2[0]\, B => 
        \wait_count_xhdl31[1]_net_1\, Y => \current_state_ns[3]\);
    
    \current_state_ns_0_a2_0[5]\ : CFG3
      generic map(INIT => x"82")

      port map(A => \current_state[2]_net_1\, B => 
        synchronizer_1_0, C => post_sync_1_reg, Y => N_359);
    
    \hwdata_r_xhdl4[9]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(9), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(9));
    
    \RD_DATA_d1[28]\ : SLE
      port map(D => rdch_read_data(28), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(28));
    
    \HADDR_d_xhdl13[19]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(19), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(19));
    
    rdch_fifo_rd_en_r_d : SLE
      port map(D => \rdch_fifo_rd_en_r\, CLK => SDRCLK_c, EN => 
        VCC_net_1, ALn => ARESET_n, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rdch_fifo_rd_en_r_d\);
    
    \current_state_RNO[7]\ : CFG4
      generic map(INIT => x"CEEE")

      port map(A => \current_state_ns_i_0_o2[1]_net_1\, B => 
        \current_state[1]_net_1\, C => masterAddrInProg_0, D => 
        N_149_i_1, Y => N_149_i);
    
    \RD_DATA_d1[7]\ : SLE
      port map(D => rdch_read_data(7), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(7));
    
    \RD_DATA_d1[18]\ : SLE
      port map(D => rdch_read_data(18), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(18));
    
    \hwdata_r_xhdl4[21]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(21), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(21));
    
    \current_state_ns_0[7]\ : CFG4
      generic map(INIT => x"FDF0")

      port map(A => \wait_count_xhdl31[1]_net_1\, B => 
        \wait_count_xhdl31[0]_net_1\, C => N_357, D => 
        \current_state[0]_net_1\, Y => \current_state_ns[7]\);
    
    ahb_busyidle_cyc_xhdl21_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \HTRANS_d_xhdl16[1]_net_1\, Y => 
        \HTRANS_d_xhdl16_i[1]\);
    
    \hwdata_r_xhdl4[19]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HWDATA(19), CLK => 
        SDRCLK_c, EN => VCC_net_1, ALn => ARESET_n, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => wrch_hwdata_r(19));
    
    \HADDR_d_xhdl13[18]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(18), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(18));
    
    \RD_DATA_d1[20]\ : SLE
      port map(D => rdch_read_data(20), CLK => SDRCLK_c, EN => 
        \rdch_fifo_rd_en_r_d\, ALn => ARESET_n, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => CoreAHBLite_0_AHBmslave10_HRDATA(20));
    
    rdch_fifo_rd_en_r_xhdl6_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => fifo_rd_en_xhdl40_1_sqmuxa, B => 
        un1_current_state_2_i, Y => N_335_i);
    
    \HADDR_d_xhdl13[0]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(0), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(0));
    
    \HSIZE_d_xhdl17[1]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HSIZE(1), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HSIZE_d(1));
    
    \HADDR_d_xhdl13[25]\ : SLE
      port map(D => CoreAHBLite_0_AHBmslave10_HADDR(25), CLK => 
        SDRCLK_c, EN => latchahbcmd_xhdl34_1, ALn => ARESET_n, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => HADDR_d(25));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI is

    port( COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : out   std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : out   std_logic_vector(27 downto 1);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : in    std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : out   std_logic_vector(63 downto 16);
          CoreAHBLite_0_AHBmslave10_HWDATA     : in    std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HRDATA     : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE      : in    std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HADDR      : in    std_logic_vector(27 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : out   std_logic;
          axi_current_state_0                  : out   std_logic;
          axi_current_state_3                  : out   std_logic;
          current_state_0                      : out   std_logic;
          masterAddrInProg_0                   : in    std_logic;
          xhdl1222_0                           : in    std_logic;
          MSS_READY                            : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : out   std_logic;
          awaddr_awvalid_clr_d                 : out   std_logic;
          araddr_arvalid_clr_d                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : in    std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : out   std_logic;
          N_75_i                               : out   std_logic;
          N_48                                 : out   std_logic;
          N_1445_i                             : out   std_logic;
          wready_m_xhdl2                       : in    std_logic;
          N_1446_i                             : out   std_logic;
          N_1452_i                             : out   std_logic;
          N_1447_i                             : out   std_logic;
          N_1451_i                             : out   std_logic;
          N_135_i                              : out   std_logic;
          N_136_i                              : out   std_logic;
          N_137_i                              : out   std_logic;
          N_203_i                              : out   std_logic;
          N_272_i                              : out   std_logic;
          N_273_i                              : out   std_logic;
          N_274_i                              : out   std_logic;
          N_275_i                              : out   std_logic;
          N_276_i                              : out   std_logic;
          N_277_i                              : out   std_logic;
          N_382_i                              : out   std_logic;
          N_381_i                              : out   std_logic;
          N_278_i                              : out   std_logic;
          N_380_i                              : out   std_logic;
          N_133_i                              : out   std_logic;
          N_134_i                              : out   std_logic;
          N_195_i                              : out   std_logic;
          N_197_i                              : out   std_logic;
          N_200_i                              : out   std_logic;
          N_201_i                              : out   std_logic;
          N_202_i                              : out   std_logic;
          N_1450_i                             : out   std_logic;
          N_1449_i                             : out   std_logic;
          N_1448_i                             : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : in    std_logic;
          SDRCLK_c                             : in    std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE     : in    std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK  : in    std_logic;
          hsel2_0_a2_1                         : in    std_logic;
          hsel2                                : in    std_logic;
          N_91                                 : in    std_logic;
          m0PrevDataSlaveReady                 : in    std_logic;
          N_92                                 : in    std_logic
        );

end top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI;

architecture DEF_ARCH of top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI is 

  component Synchronizer_AHBtoAXIHX
    port( N_163_i            : in    std_logic := 'U';
          ahb_rd_req_sync    : out   std_logic;
          latch_ahb_sig      : in    std_logic := 'U';
          latch_ahb_sig_sync : out   std_logic;
          ahb_wr_done        : in    std_logic := 'U';
          wrch_fifo_wr_en_r  : out   std_logic;
          SDRCLK_c           : in    std_logic := 'U';
          ARESET_n           : in    std_logic := 'U';
          ahb_wr_done_sync   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CoreAHBLtoAXI_WRCHANNELFIFOHX
    port( wrch_hwdata_r       : in    std_logic_vector(31 downto 0) := (others => 'U');
          masterAddrInProg_0  : in    std_logic := 'U';
          axi_current_state_0 : in    std_logic := 'U';
          valid_ahbcmd_i_o3_1 : in    std_logic := 'U';
          hsel2_0_a2_1        : in    std_logic := 'U';
          N_209               : out   std_logic;
          N_210               : out   std_logic;
          N_213               : out   std_logic;
          N_214               : out   std_logic;
          N_215               : out   std_logic;
          N_217               : out   std_logic;
          N_218               : out   std_logic;
          N_221               : out   std_logic;
          N_222               : out   std_logic;
          N_223               : out   std_logic;
          N_328               : out   std_logic;
          N_440               : out   std_logic;
          N_439               : out   std_logic;
          N_438               : out   std_logic;
          N_437               : out   std_logic;
          N_436               : out   std_logic;
          N_435               : out   std_logic;
          N_434               : out   std_logic;
          N_433               : out   std_logic;
          N_432               : out   std_logic;
          N_431               : out   std_logic;
          N_430               : out   std_logic;
          N_429               : out   std_logic;
          N_428               : out   std_logic;
          N_427               : out   std_logic;
          N_426               : out   std_logic;
          N_425               : out   std_logic;
          N_424               : out   std_logic;
          N_423               : out   std_logic;
          N_422               : out   std_logic;
          N_421               : out   std_logic;
          N_420               : out   std_logic;
          N_419               : out   std_logic;
          N_418               : out   std_logic;
          N_417               : out   std_logic;
          N_416               : out   std_logic;
          N_415               : out   std_logic;
          N_414               : out   std_logic;
          N_413               : out   std_logic;
          N_412               : out   std_logic;
          N_411               : out   std_logic;
          N_410               : out   std_logic;
          N_293               : out   std_logic;
          N_292               : out   std_logic;
          N_291               : out   std_logic;
          N_290               : out   std_logic;
          N_289               : out   std_logic;
          N_288               : out   std_logic;
          N_286               : out   std_logic;
          N_285               : out   std_logic;
          N_284               : out   std_logic;
          N_283               : out   std_logic;
          N_282               : out   std_logic;
          N_281               : out   std_logic;
          N_160               : out   std_logic;
          N_159               : out   std_logic;
          N_158               : out   std_logic;
          N_157               : out   std_logic;
          N_156               : out   std_logic;
          N_151               : out   std_logic;
          N_150               : out   std_logic;
          N_149               : out   std_logic;
          N_148               : out   std_logic;
          N_147               : out   std_logic;
          wrch_fifo_wr_en_r   : in    std_logic := 'U';
          ahb_busyidle_cyc    : in    std_logic := 'U';
          N_72_i              : in    std_logic := 'U';
          N_98                : in    std_logic := 'U';
          N_73_i_0            : in    std_logic := 'U';
          ahb_busyidle_cyc_i  : in    std_logic := 'U';
          SDRCLK_c            : in    std_logic := 'U';
          ARESET_n            : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLtoAXI_reset_syncHX_0
    port( SDRCLK_c  : in    std_logic := 'U';
          MSS_READY : in    std_logic := 'U';
          ARESET_n  : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CoreAHBLtoAXI_RDCHANNELFIFOHX
    port( rdch_read_data      : out   std_logic_vector(31 downto 0);
          rdch_fifo_wr_data   : in    std_logic_vector(31 downto 0) := (others => 'U');
          masterAddrInProg_0  : in    std_logic := 'U';
          valid_ahbcmd_i_o3_1 : in    std_logic := 'U';
          hsel2_0_a2_1        : in    std_logic := 'U';
          rdch_fifo_wr_en_r   : in    std_logic := 'U';
          rdch_fifo_rd_en_r   : in    std_logic := 'U';
          rdch_fifo_empty     : out   std_logic;
          SDRCLK_c            : in    std_logic := 'U';
          ARESET_n            : in    std_logic := 'U'
        );
  end component;

  component Synchronizer_AXItoAHBHX
    port( synchronizer_1_0                   : out   std_logic;
          BVALID_sync                        : out   std_logic;
          axi_read_rlast                     : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_BVALID : in    std_logic := 'U';
          post_sync_1_reg                    : out   std_logic;
          SDRCLK_c                           : in    std_logic := 'U';
          ARESET_n                           : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLtoAXI_AXIAccessControlHX
    port( COREAHBLTOAXI_0_AXIMasterIF_WDATA    : out   std_logic_vector(63 downto 16);
          rdch_fifo_wr_data                    : out   std_logic_vector(31 downto 0);
          HADDR_d                              : in    std_logic_vector(27 downto 0) := (others => 'U');
          HSIZE_d                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : in    std_logic_vector(63 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : out   std_logic_vector(27 downto 1);
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : out   std_logic_vector(1 downto 0);
          axi_current_state_0                  : out   std_logic;
          axi_current_state_3                  : out   std_logic;
          axi_current_state_2                  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : out   std_logic;
          N_1448_i                             : out   std_logic;
          N_1449_i                             : out   std_logic;
          N_1450_i                             : out   std_logic;
          N_202_i                              : out   std_logic;
          N_201_i                              : out   std_logic;
          N_200_i                              : out   std_logic;
          N_197_i                              : out   std_logic;
          N_195_i                              : out   std_logic;
          N_134_i                              : out   std_logic;
          N_133_i                              : out   std_logic;
          N_380_i                              : out   std_logic;
          N_278_i                              : out   std_logic;
          N_381_i                              : out   std_logic;
          N_382_i                              : out   std_logic;
          N_277_i                              : out   std_logic;
          N_276_i                              : out   std_logic;
          N_275_i                              : out   std_logic;
          N_274_i                              : out   std_logic;
          N_273_i                              : out   std_logic;
          N_272_i                              : out   std_logic;
          N_203_i                              : out   std_logic;
          N_137_i                              : out   std_logic;
          N_136_i                              : out   std_logic;
          N_135_i                              : out   std_logic;
          N_209                                : in    std_logic := 'U';
          N_217                                : in    std_logic := 'U';
          N_210                                : in    std_logic := 'U';
          N_218                                : in    std_logic := 'U';
          N_213                                : in    std_logic := 'U';
          N_221                                : in    std_logic := 'U';
          N_214                                : in    std_logic := 'U';
          N_222                                : in    std_logic := 'U';
          N_215                                : in    std_logic := 'U';
          N_223                                : in    std_logic := 'U';
          N_432                                : in    std_logic := 'U';
          N_439                                : in    std_logic := 'U';
          N_431                                : in    std_logic := 'U';
          N_438                                : in    std_logic := 'U';
          N_430                                : in    std_logic := 'U';
          N_437                                : in    std_logic := 'U';
          N_429                                : in    std_logic := 'U';
          N_436                                : in    std_logic := 'U';
          N_428                                : in    std_logic := 'U';
          N_435                                : in    std_logic := 'U';
          N_427                                : in    std_logic := 'U';
          N_434                                : in    std_logic := 'U';
          N_426                                : in    std_logic := 'U';
          N_433                                : in    std_logic := 'U';
          N_421                                : in    std_logic := 'U';
          N_425                                : in    std_logic := 'U';
          N_420                                : in    std_logic := 'U';
          N_424                                : in    std_logic := 'U';
          N_419                                : in    std_logic := 'U';
          N_423                                : in    std_logic := 'U';
          N_418                                : in    std_logic := 'U';
          N_422                                : in    std_logic := 'U';
          N_417                                : in    std_logic := 'U';
          N_414                                : in    std_logic := 'U';
          N_416                                : in    std_logic := 'U';
          N_413                                : in    std_logic := 'U';
          N_328                                : in    std_logic := 'U';
          N_440                                : in    std_logic := 'U';
          N_412                                : in    std_logic := 'U';
          N_415                                : in    std_logic := 'U';
          N_410                                : in    std_logic := 'U';
          N_411                                : in    std_logic := 'U';
          N_286                                : in    std_logic := 'U';
          N_293                                : in    std_logic := 'U';
          N_285                                : in    std_logic := 'U';
          N_292                                : in    std_logic := 'U';
          N_284                                : in    std_logic := 'U';
          N_291                                : in    std_logic := 'U';
          N_283                                : in    std_logic := 'U';
          N_290                                : in    std_logic := 'U';
          N_282                                : in    std_logic := 'U';
          N_289                                : in    std_logic := 'U';
          N_281                                : in    std_logic := 'U';
          N_288                                : in    std_logic := 'U';
          N_151                                : in    std_logic := 'U';
          N_160                                : in    std_logic := 'U';
          N_150                                : in    std_logic := 'U';
          N_159                                : in    std_logic := 'U';
          N_149                                : in    std_logic := 'U';
          N_158                                : in    std_logic := 'U';
          N_148                                : in    std_logic := 'U';
          N_157                                : in    std_logic := 'U';
          N_147                                : in    std_logic := 'U';
          N_156                                : in    std_logic := 'U';
          N_1451_i                             : out   std_logic;
          N_1447_i                             : out   std_logic;
          N_1452_i                             : out   std_logic;
          N_1446_i                             : out   std_logic;
          wready_m_xhdl2                       : in    std_logic := 'U';
          N_73_i_0                             : out   std_logic;
          N_72_i                               : out   std_logic;
          N_1445_i                             : out   std_logic;
          N_48                                 : out   std_logic;
          N_75_i                               : out   std_logic;
          ahb_wr_done_sync                     : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic := 'U';
          N_98                                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : in    std_logic := 'U';
          araddr_arvalid_clr_d                 : out   std_logic;
          awaddr_awvalid_clr_d                 : out   std_logic;
          ahb_rd_req_sync                      : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : in    std_logic := 'U';
          latch_ahb_sig_sync                   : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : out   std_logic;
          rdch_fifo_wr_en_r                    : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : out   std_logic;
          axi_read_rlast                       : out   std_logic;
          HMASTLOCK_d                          : in    std_logic := 'U';
          HWRITE_d                             : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          ARESET_n                             : in    std_logic := 'U'
        );
  end component;

  component CoreAHBLtoAXI_AHBAccessControlHX
    port( CoreAHBLite_0_AHBmslave10_HADDR     : in    std_logic_vector(27 downto 0) := (others => 'U');
          HADDR_d                             : out   std_logic_vector(27 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE     : in    std_logic_vector(1 downto 0) := (others => 'U');
          HSIZE_d                             : out   std_logic_vector(1 downto 0);
          rdch_read_data                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HRDATA    : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA    : in    std_logic_vector(31 downto 0) := (others => 'U');
          wrch_hwdata_r                       : out   std_logic_vector(31 downto 0);
          xhdl1222_0                          : in    std_logic := 'U';
          synchronizer_1_0                    : in    std_logic := 'U';
          masterAddrInProg_0                  : in    std_logic := 'U';
          current_state_0                     : out   std_logic;
          N_92                                : in    std_logic := 'U';
          m0PrevDataSlaveReady                : in    std_logic := 'U';
          N_91                                : in    std_logic := 'U';
          post_sync_1_reg                     : in    std_logic := 'U';
          rdch_fifo_empty                     : in    std_logic := 'U';
          N_163_i                             : out   std_logic;
          hsel2                               : in    std_logic := 'U';
          hsel2_0_a2_1                        : in    std_logic := 'U';
          valid_ahbcmd_i_o3_1                 : out   std_logic;
          rdch_fifo_rd_en_r                   : out   std_logic;
          latch_ahb_sig                       : out   std_logic;
          BVALID_sync                         : in    std_logic := 'U';
          ahb_wr_done                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HMASTLOCK : in    std_logic := 'U';
          HMASTLOCK_d                         : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE    : in    std_logic := 'U';
          HWRITE_d                            : out   std_logic;
          SDRCLK_c                            : in    std_logic := 'U';
          ARESET_n                            : in    std_logic := 'U';
          ahb_busyidle_cyc_i                  : out   std_logic;
          ahb_busyidle_cyc                    : out   std_logic
        );
  end component;

    signal \synchronizer_1[0]\, \HADDR_d[0]\, \HADDR_d[1]\, 
        \HADDR_d[2]\, \HADDR_d[3]\, \HADDR_d[4]\, \HADDR_d[5]\, 
        \HADDR_d[6]\, \HADDR_d[7]\, \HADDR_d[8]\, \HADDR_d[9]\, 
        \HADDR_d[10]\, \HADDR_d[11]\, \HADDR_d[12]\, 
        \HADDR_d[13]\, \HADDR_d[14]\, \HADDR_d[15]\, 
        \HADDR_d[16]\, \HADDR_d[17]\, \HADDR_d[18]\, 
        \HADDR_d[19]\, \HADDR_d[20]\, \HADDR_d[21]\, 
        \HADDR_d[22]\, \HADDR_d[23]\, \HADDR_d[24]\, 
        \HADDR_d[25]\, \HADDR_d[26]\, \HADDR_d[27]\, \HSIZE_d[0]\, 
        \HSIZE_d[1]\, \rdch_read_data[0]\, \rdch_read_data[1]\, 
        \rdch_read_data[2]\, \rdch_read_data[3]\, 
        \rdch_read_data[4]\, \rdch_read_data[5]\, 
        \rdch_read_data[6]\, \rdch_read_data[7]\, 
        \rdch_read_data[8]\, \rdch_read_data[9]\, 
        \rdch_read_data[10]\, \rdch_read_data[11]\, 
        \rdch_read_data[12]\, \rdch_read_data[13]\, 
        \rdch_read_data[14]\, \rdch_read_data[15]\, 
        \rdch_read_data[16]\, \rdch_read_data[17]\, 
        \rdch_read_data[18]\, \rdch_read_data[19]\, 
        \rdch_read_data[20]\, \rdch_read_data[21]\, 
        \rdch_read_data[22]\, \rdch_read_data[23]\, 
        \rdch_read_data[24]\, \rdch_read_data[25]\, 
        \rdch_read_data[26]\, \rdch_read_data[27]\, 
        \rdch_read_data[28]\, \rdch_read_data[29]\, 
        \rdch_read_data[30]\, \rdch_read_data[31]\, 
        \wrch_hwdata_r[0]\, \wrch_hwdata_r[1]\, 
        \wrch_hwdata_r[2]\, \wrch_hwdata_r[3]\, 
        \wrch_hwdata_r[4]\, \wrch_hwdata_r[5]\, 
        \wrch_hwdata_r[6]\, \wrch_hwdata_r[7]\, 
        \wrch_hwdata_r[8]\, \wrch_hwdata_r[9]\, 
        \wrch_hwdata_r[10]\, \wrch_hwdata_r[11]\, 
        \wrch_hwdata_r[12]\, \wrch_hwdata_r[13]\, 
        \wrch_hwdata_r[14]\, \wrch_hwdata_r[15]\, 
        \wrch_hwdata_r[16]\, \wrch_hwdata_r[17]\, 
        \wrch_hwdata_r[18]\, \wrch_hwdata_r[19]\, 
        \wrch_hwdata_r[20]\, \wrch_hwdata_r[21]\, 
        \wrch_hwdata_r[22]\, \wrch_hwdata_r[23]\, 
        \wrch_hwdata_r[24]\, \wrch_hwdata_r[25]\, 
        \wrch_hwdata_r[26]\, \wrch_hwdata_r[27]\, 
        \wrch_hwdata_r[28]\, \wrch_hwdata_r[29]\, 
        \wrch_hwdata_r[30]\, \wrch_hwdata_r[31]\, post_sync_1_reg, 
        rdch_fifo_empty, N_163_i, valid_ahbcmd_i_o3_1, 
        rdch_fifo_rd_en_r, latch_ahb_sig, BVALID_sync, 
        ahb_wr_done, HMASTLOCK_d, HWRITE_d, ARESET_n, 
        ahb_busyidle_cyc_i, ahb_busyidle_cyc, 
        \axi_current_state[3]\, N_209, N_210, N_213, N_214, N_215, 
        N_217, N_218, N_221, N_222, N_223, N_328, N_440, N_439, 
        N_438, N_437, N_436, N_435, N_434, N_433, N_432, N_431, 
        N_430, N_429, N_428, N_427, N_426, N_425, N_424, N_423, 
        N_422, N_421, N_420, N_419, N_418, N_417, N_416, N_415, 
        N_414, N_413, N_412, N_411, N_410, N_293, N_292, N_291, 
        N_290, N_289, N_288, N_286, N_285, N_284, N_283, N_282, 
        N_281, N_160, N_159, N_158, N_157, N_156, N_151, N_150, 
        N_149, N_148, N_147, wrch_fifo_wr_en_r, N_72_i, N_98, 
        N_73_i_0, ahb_rd_req_sync, latch_ahb_sig_sync, 
        ahb_wr_done_sync, axi_read_rlast, \rdch_fifo_wr_data[0]\, 
        \rdch_fifo_wr_data[1]\, \rdch_fifo_wr_data[2]\, 
        \rdch_fifo_wr_data[3]\, \rdch_fifo_wr_data[4]\, 
        \rdch_fifo_wr_data[5]\, \rdch_fifo_wr_data[6]\, 
        \rdch_fifo_wr_data[7]\, \rdch_fifo_wr_data[8]\, 
        \rdch_fifo_wr_data[9]\, \rdch_fifo_wr_data[10]\, 
        \rdch_fifo_wr_data[11]\, \rdch_fifo_wr_data[12]\, 
        \rdch_fifo_wr_data[13]\, \rdch_fifo_wr_data[14]\, 
        \rdch_fifo_wr_data[15]\, \rdch_fifo_wr_data[16]\, 
        \rdch_fifo_wr_data[17]\, \rdch_fifo_wr_data[18]\, 
        \rdch_fifo_wr_data[19]\, \rdch_fifo_wr_data[20]\, 
        \rdch_fifo_wr_data[21]\, \rdch_fifo_wr_data[22]\, 
        \rdch_fifo_wr_data[23]\, \rdch_fifo_wr_data[24]\, 
        \rdch_fifo_wr_data[25]\, \rdch_fifo_wr_data[26]\, 
        \rdch_fifo_wr_data[27]\, \rdch_fifo_wr_data[28]\, 
        \rdch_fifo_wr_data[29]\, \rdch_fifo_wr_data[30]\, 
        \rdch_fifo_wr_data[31]\, rdch_fifo_wr_en_r, GND_net_1, 
        VCC_net_1 : std_logic;
    signal nc2, nc5, nc4, nc3, nc1 : std_logic;

    for all : Synchronizer_AHBtoAXIHX
	Use entity work.Synchronizer_AHBtoAXIHX(DEF_ARCH);
    for all : CoreAHBLtoAXI_WRCHANNELFIFOHX
	Use entity work.CoreAHBLtoAXI_WRCHANNELFIFOHX(DEF_ARCH);
    for all : CoreAHBLtoAXI_reset_syncHX_0
	Use entity work.CoreAHBLtoAXI_reset_syncHX_0(DEF_ARCH);
    for all : CoreAHBLtoAXI_RDCHANNELFIFOHX
	Use entity work.CoreAHBLtoAXI_RDCHANNELFIFOHX(DEF_ARCH);
    for all : Synchronizer_AXItoAHBHX
	Use entity work.Synchronizer_AXItoAHBHX(DEF_ARCH);
    for all : CoreAHBLtoAXI_AXIAccessControlHX
	Use entity work.CoreAHBLtoAXI_AXIAccessControlHX(DEF_ARCH);
    for all : CoreAHBLtoAXI_AHBAccessControlHX
	Use entity work.CoreAHBLtoAXI_AHBAccessControlHX(DEF_ARCH);
begin 


    U_AHBtoAXI_sync : Synchronizer_AHBtoAXIHX
      port map(N_163_i => N_163_i, ahb_rd_req_sync => 
        ahb_rd_req_sync, latch_ahb_sig => latch_ahb_sig, 
        latch_ahb_sig_sync => latch_ahb_sig_sync, ahb_wr_done => 
        ahb_wr_done, wrch_fifo_wr_en_r => wrch_fifo_wr_en_r, 
        SDRCLK_c => SDRCLK_c, ARESET_n => ARESET_n, 
        ahb_wr_done_sync => ahb_wr_done_sync);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U_WrChannelFifo : CoreAHBLtoAXI_WRCHANNELFIFOHX
      port map(wrch_hwdata_r(31) => \wrch_hwdata_r[31]\, 
        wrch_hwdata_r(30) => \wrch_hwdata_r[30]\, 
        wrch_hwdata_r(29) => \wrch_hwdata_r[29]\, 
        wrch_hwdata_r(28) => \wrch_hwdata_r[28]\, 
        wrch_hwdata_r(27) => \wrch_hwdata_r[27]\, 
        wrch_hwdata_r(26) => \wrch_hwdata_r[26]\, 
        wrch_hwdata_r(25) => \wrch_hwdata_r[25]\, 
        wrch_hwdata_r(24) => \wrch_hwdata_r[24]\, 
        wrch_hwdata_r(23) => \wrch_hwdata_r[23]\, 
        wrch_hwdata_r(22) => \wrch_hwdata_r[22]\, 
        wrch_hwdata_r(21) => \wrch_hwdata_r[21]\, 
        wrch_hwdata_r(20) => \wrch_hwdata_r[20]\, 
        wrch_hwdata_r(19) => \wrch_hwdata_r[19]\, 
        wrch_hwdata_r(18) => \wrch_hwdata_r[18]\, 
        wrch_hwdata_r(17) => \wrch_hwdata_r[17]\, 
        wrch_hwdata_r(16) => \wrch_hwdata_r[16]\, 
        wrch_hwdata_r(15) => \wrch_hwdata_r[15]\, 
        wrch_hwdata_r(14) => \wrch_hwdata_r[14]\, 
        wrch_hwdata_r(13) => \wrch_hwdata_r[13]\, 
        wrch_hwdata_r(12) => \wrch_hwdata_r[12]\, 
        wrch_hwdata_r(11) => \wrch_hwdata_r[11]\, 
        wrch_hwdata_r(10) => \wrch_hwdata_r[10]\, 
        wrch_hwdata_r(9) => \wrch_hwdata_r[9]\, wrch_hwdata_r(8)
         => \wrch_hwdata_r[8]\, wrch_hwdata_r(7) => 
        \wrch_hwdata_r[7]\, wrch_hwdata_r(6) => 
        \wrch_hwdata_r[6]\, wrch_hwdata_r(5) => 
        \wrch_hwdata_r[5]\, wrch_hwdata_r(4) => 
        \wrch_hwdata_r[4]\, wrch_hwdata_r(3) => 
        \wrch_hwdata_r[3]\, wrch_hwdata_r(2) => 
        \wrch_hwdata_r[2]\, wrch_hwdata_r(1) => 
        \wrch_hwdata_r[1]\, wrch_hwdata_r(0) => 
        \wrch_hwdata_r[0]\, masterAddrInProg_0 => 
        masterAddrInProg_0, axi_current_state_0 => 
        \axi_current_state[3]\, valid_ahbcmd_i_o3_1 => 
        valid_ahbcmd_i_o3_1, hsel2_0_a2_1 => hsel2_0_a2_1, N_209
         => N_209, N_210 => N_210, N_213 => N_213, N_214 => N_214, 
        N_215 => N_215, N_217 => N_217, N_218 => N_218, N_221 => 
        N_221, N_222 => N_222, N_223 => N_223, N_328 => N_328, 
        N_440 => N_440, N_439 => N_439, N_438 => N_438, N_437 => 
        N_437, N_436 => N_436, N_435 => N_435, N_434 => N_434, 
        N_433 => N_433, N_432 => N_432, N_431 => N_431, N_430 => 
        N_430, N_429 => N_429, N_428 => N_428, N_427 => N_427, 
        N_426 => N_426, N_425 => N_425, N_424 => N_424, N_423 => 
        N_423, N_422 => N_422, N_421 => N_421, N_420 => N_420, 
        N_419 => N_419, N_418 => N_418, N_417 => N_417, N_416 => 
        N_416, N_415 => N_415, N_414 => N_414, N_413 => N_413, 
        N_412 => N_412, N_411 => N_411, N_410 => N_410, N_293 => 
        N_293, N_292 => N_292, N_291 => N_291, N_290 => N_290, 
        N_289 => N_289, N_288 => N_288, N_286 => N_286, N_285 => 
        N_285, N_284 => N_284, N_283 => N_283, N_282 => N_282, 
        N_281 => N_281, N_160 => N_160, N_159 => N_159, N_158 => 
        N_158, N_157 => N_157, N_156 => N_156, N_151 => N_151, 
        N_150 => N_150, N_149 => N_149, N_148 => N_148, N_147 => 
        N_147, wrch_fifo_wr_en_r => wrch_fifo_wr_en_r, 
        ahb_busyidle_cyc => ahb_busyidle_cyc, N_72_i => N_72_i, 
        N_98 => N_98, N_73_i_0 => N_73_i_0, ahb_busyidle_cyc_i
         => ahb_busyidle_cyc_i, SDRCLK_c => SDRCLK_c, ARESET_n
         => ARESET_n);
    
    U_RST_A : CoreAHBLtoAXI_reset_syncHX_0
      port map(SDRCLK_c => SDRCLK_c, MSS_READY => MSS_READY, 
        ARESET_n => ARESET_n);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U_RdChannelFifo : CoreAHBLtoAXI_RDCHANNELFIFOHX
      port map(rdch_read_data(31) => \rdch_read_data[31]\, 
        rdch_read_data(30) => \rdch_read_data[30]\, 
        rdch_read_data(29) => \rdch_read_data[29]\, 
        rdch_read_data(28) => \rdch_read_data[28]\, 
        rdch_read_data(27) => \rdch_read_data[27]\, 
        rdch_read_data(26) => \rdch_read_data[26]\, 
        rdch_read_data(25) => \rdch_read_data[25]\, 
        rdch_read_data(24) => \rdch_read_data[24]\, 
        rdch_read_data(23) => \rdch_read_data[23]\, 
        rdch_read_data(22) => \rdch_read_data[22]\, 
        rdch_read_data(21) => \rdch_read_data[21]\, 
        rdch_read_data(20) => \rdch_read_data[20]\, 
        rdch_read_data(19) => \rdch_read_data[19]\, 
        rdch_read_data(18) => \rdch_read_data[18]\, 
        rdch_read_data(17) => \rdch_read_data[17]\, 
        rdch_read_data(16) => \rdch_read_data[16]\, 
        rdch_read_data(15) => \rdch_read_data[15]\, 
        rdch_read_data(14) => \rdch_read_data[14]\, 
        rdch_read_data(13) => \rdch_read_data[13]\, 
        rdch_read_data(12) => \rdch_read_data[12]\, 
        rdch_read_data(11) => \rdch_read_data[11]\, 
        rdch_read_data(10) => \rdch_read_data[10]\, 
        rdch_read_data(9) => \rdch_read_data[9]\, 
        rdch_read_data(8) => \rdch_read_data[8]\, 
        rdch_read_data(7) => \rdch_read_data[7]\, 
        rdch_read_data(6) => \rdch_read_data[6]\, 
        rdch_read_data(5) => \rdch_read_data[5]\, 
        rdch_read_data(4) => \rdch_read_data[4]\, 
        rdch_read_data(3) => \rdch_read_data[3]\, 
        rdch_read_data(2) => \rdch_read_data[2]\, 
        rdch_read_data(1) => \rdch_read_data[1]\, 
        rdch_read_data(0) => \rdch_read_data[0]\, 
        rdch_fifo_wr_data(31) => \rdch_fifo_wr_data[31]\, 
        rdch_fifo_wr_data(30) => \rdch_fifo_wr_data[30]\, 
        rdch_fifo_wr_data(29) => \rdch_fifo_wr_data[29]\, 
        rdch_fifo_wr_data(28) => \rdch_fifo_wr_data[28]\, 
        rdch_fifo_wr_data(27) => \rdch_fifo_wr_data[27]\, 
        rdch_fifo_wr_data(26) => \rdch_fifo_wr_data[26]\, 
        rdch_fifo_wr_data(25) => \rdch_fifo_wr_data[25]\, 
        rdch_fifo_wr_data(24) => \rdch_fifo_wr_data[24]\, 
        rdch_fifo_wr_data(23) => \rdch_fifo_wr_data[23]\, 
        rdch_fifo_wr_data(22) => \rdch_fifo_wr_data[22]\, 
        rdch_fifo_wr_data(21) => \rdch_fifo_wr_data[21]\, 
        rdch_fifo_wr_data(20) => \rdch_fifo_wr_data[20]\, 
        rdch_fifo_wr_data(19) => \rdch_fifo_wr_data[19]\, 
        rdch_fifo_wr_data(18) => \rdch_fifo_wr_data[18]\, 
        rdch_fifo_wr_data(17) => \rdch_fifo_wr_data[17]\, 
        rdch_fifo_wr_data(16) => \rdch_fifo_wr_data[16]\, 
        rdch_fifo_wr_data(15) => \rdch_fifo_wr_data[15]\, 
        rdch_fifo_wr_data(14) => \rdch_fifo_wr_data[14]\, 
        rdch_fifo_wr_data(13) => \rdch_fifo_wr_data[13]\, 
        rdch_fifo_wr_data(12) => \rdch_fifo_wr_data[12]\, 
        rdch_fifo_wr_data(11) => \rdch_fifo_wr_data[11]\, 
        rdch_fifo_wr_data(10) => \rdch_fifo_wr_data[10]\, 
        rdch_fifo_wr_data(9) => \rdch_fifo_wr_data[9]\, 
        rdch_fifo_wr_data(8) => \rdch_fifo_wr_data[8]\, 
        rdch_fifo_wr_data(7) => \rdch_fifo_wr_data[7]\, 
        rdch_fifo_wr_data(6) => \rdch_fifo_wr_data[6]\, 
        rdch_fifo_wr_data(5) => \rdch_fifo_wr_data[5]\, 
        rdch_fifo_wr_data(4) => \rdch_fifo_wr_data[4]\, 
        rdch_fifo_wr_data(3) => \rdch_fifo_wr_data[3]\, 
        rdch_fifo_wr_data(2) => \rdch_fifo_wr_data[2]\, 
        rdch_fifo_wr_data(1) => \rdch_fifo_wr_data[1]\, 
        rdch_fifo_wr_data(0) => \rdch_fifo_wr_data[0]\, 
        masterAddrInProg_0 => masterAddrInProg_0, 
        valid_ahbcmd_i_o3_1 => valid_ahbcmd_i_o3_1, hsel2_0_a2_1
         => hsel2_0_a2_1, rdch_fifo_wr_en_r => rdch_fifo_wr_en_r, 
        rdch_fifo_rd_en_r => rdch_fifo_rd_en_r, rdch_fifo_empty
         => rdch_fifo_empty, SDRCLK_c => SDRCLK_c, ARESET_n => 
        ARESET_n);
    
    U_AXItoAHB_sync : Synchronizer_AXItoAHBHX
      port map(synchronizer_1_0 => \synchronizer_1[0]\, 
        BVALID_sync => BVALID_sync, axi_read_rlast => 
        axi_read_rlast, COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID, post_sync_1_reg => 
        post_sync_1_reg, SDRCLK_c => SDRCLK_c, ARESET_n => 
        ARESET_n);
    
    U_AXIAccCntrl : CoreAHBLtoAXI_AXIAccessControlHX
      port map(COREAHBLTOAXI_0_AXIMasterIF_WDATA(63) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(63), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(31) => nc2, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(28) => nc5, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(21) => nc4, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(20) => nc3, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(19) => nc1, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17), 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16), 
        rdch_fifo_wr_data(31) => \rdch_fifo_wr_data[31]\, 
        rdch_fifo_wr_data(30) => \rdch_fifo_wr_data[30]\, 
        rdch_fifo_wr_data(29) => \rdch_fifo_wr_data[29]\, 
        rdch_fifo_wr_data(28) => \rdch_fifo_wr_data[28]\, 
        rdch_fifo_wr_data(27) => \rdch_fifo_wr_data[27]\, 
        rdch_fifo_wr_data(26) => \rdch_fifo_wr_data[26]\, 
        rdch_fifo_wr_data(25) => \rdch_fifo_wr_data[25]\, 
        rdch_fifo_wr_data(24) => \rdch_fifo_wr_data[24]\, 
        rdch_fifo_wr_data(23) => \rdch_fifo_wr_data[23]\, 
        rdch_fifo_wr_data(22) => \rdch_fifo_wr_data[22]\, 
        rdch_fifo_wr_data(21) => \rdch_fifo_wr_data[21]\, 
        rdch_fifo_wr_data(20) => \rdch_fifo_wr_data[20]\, 
        rdch_fifo_wr_data(19) => \rdch_fifo_wr_data[19]\, 
        rdch_fifo_wr_data(18) => \rdch_fifo_wr_data[18]\, 
        rdch_fifo_wr_data(17) => \rdch_fifo_wr_data[17]\, 
        rdch_fifo_wr_data(16) => \rdch_fifo_wr_data[16]\, 
        rdch_fifo_wr_data(15) => \rdch_fifo_wr_data[15]\, 
        rdch_fifo_wr_data(14) => \rdch_fifo_wr_data[14]\, 
        rdch_fifo_wr_data(13) => \rdch_fifo_wr_data[13]\, 
        rdch_fifo_wr_data(12) => \rdch_fifo_wr_data[12]\, 
        rdch_fifo_wr_data(11) => \rdch_fifo_wr_data[11]\, 
        rdch_fifo_wr_data(10) => \rdch_fifo_wr_data[10]\, 
        rdch_fifo_wr_data(9) => \rdch_fifo_wr_data[9]\, 
        rdch_fifo_wr_data(8) => \rdch_fifo_wr_data[8]\, 
        rdch_fifo_wr_data(7) => \rdch_fifo_wr_data[7]\, 
        rdch_fifo_wr_data(6) => \rdch_fifo_wr_data[6]\, 
        rdch_fifo_wr_data(5) => \rdch_fifo_wr_data[5]\, 
        rdch_fifo_wr_data(4) => \rdch_fifo_wr_data[4]\, 
        rdch_fifo_wr_data(3) => \rdch_fifo_wr_data[3]\, 
        rdch_fifo_wr_data(2) => \rdch_fifo_wr_data[2]\, 
        rdch_fifo_wr_data(1) => \rdch_fifo_wr_data[1]\, 
        rdch_fifo_wr_data(0) => \rdch_fifo_wr_data[0]\, 
        HADDR_d(27) => \HADDR_d[27]\, HADDR_d(26) => 
        \HADDR_d[26]\, HADDR_d(25) => \HADDR_d[25]\, HADDR_d(24)
         => \HADDR_d[24]\, HADDR_d(23) => \HADDR_d[23]\, 
        HADDR_d(22) => \HADDR_d[22]\, HADDR_d(21) => 
        \HADDR_d[21]\, HADDR_d(20) => \HADDR_d[20]\, HADDR_d(19)
         => \HADDR_d[19]\, HADDR_d(18) => \HADDR_d[18]\, 
        HADDR_d(17) => \HADDR_d[17]\, HADDR_d(16) => 
        \HADDR_d[16]\, HADDR_d(15) => \HADDR_d[15]\, HADDR_d(14)
         => \HADDR_d[14]\, HADDR_d(13) => \HADDR_d[13]\, 
        HADDR_d(12) => \HADDR_d[12]\, HADDR_d(11) => 
        \HADDR_d[11]\, HADDR_d(10) => \HADDR_d[10]\, HADDR_d(9)
         => \HADDR_d[9]\, HADDR_d(8) => \HADDR_d[8]\, HADDR_d(7)
         => \HADDR_d[7]\, HADDR_d(6) => \HADDR_d[6]\, HADDR_d(5)
         => \HADDR_d[5]\, HADDR_d(4) => \HADDR_d[4]\, HADDR_d(3)
         => \HADDR_d[3]\, HADDR_d(2) => \HADDR_d[2]\, HADDR_d(1)
         => \HADDR_d[1]\, HADDR_d(0) => \HADDR_d[0]\, HSIZE_d(1)
         => \HSIZE_d[1]\, HSIZE_d(0) => \HSIZE_d[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1), 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0) => 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2), 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1), 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1), 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0) => 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0), 
        axi_current_state_0 => axi_current_state_0, 
        axi_current_state_3 => axi_current_state_3, 
        axi_current_state_2 => \axi_current_state[3]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0, N_1448_i => 
        N_1448_i, N_1449_i => N_1449_i, N_1450_i => N_1450_i, 
        N_202_i => N_202_i, N_201_i => N_201_i, N_200_i => 
        N_200_i, N_197_i => N_197_i, N_195_i => N_195_i, N_134_i
         => N_134_i, N_133_i => N_133_i, N_380_i => N_380_i, 
        N_278_i => N_278_i, N_381_i => N_381_i, N_382_i => 
        N_382_i, N_277_i => N_277_i, N_276_i => N_276_i, N_275_i
         => N_275_i, N_274_i => N_274_i, N_273_i => N_273_i, 
        N_272_i => N_272_i, N_203_i => N_203_i, N_137_i => 
        N_137_i, N_136_i => N_136_i, N_135_i => N_135_i, N_209
         => N_209, N_217 => N_217, N_210 => N_210, N_218 => N_218, 
        N_213 => N_213, N_221 => N_221, N_214 => N_214, N_222 => 
        N_222, N_215 => N_215, N_223 => N_223, N_432 => N_432, 
        N_439 => N_439, N_431 => N_431, N_438 => N_438, N_430 => 
        N_430, N_437 => N_437, N_429 => N_429, N_436 => N_436, 
        N_428 => N_428, N_435 => N_435, N_427 => N_427, N_434 => 
        N_434, N_426 => N_426, N_433 => N_433, N_421 => N_421, 
        N_425 => N_425, N_420 => N_420, N_424 => N_424, N_419 => 
        N_419, N_423 => N_423, N_418 => N_418, N_422 => N_422, 
        N_417 => N_417, N_414 => N_414, N_416 => N_416, N_413 => 
        N_413, N_328 => N_328, N_440 => N_440, N_412 => N_412, 
        N_415 => N_415, N_410 => N_410, N_411 => N_411, N_286 => 
        N_286, N_293 => N_293, N_285 => N_285, N_292 => N_292, 
        N_284 => N_284, N_291 => N_291, N_283 => N_283, N_290 => 
        N_290, N_282 => N_282, N_289 => N_289, N_281 => N_281, 
        N_288 => N_288, N_151 => N_151, N_160 => N_160, N_150 => 
        N_150, N_159 => N_159, N_149 => N_149, N_158 => N_158, 
        N_148 => N_148, N_157 => N_157, N_147 => N_147, N_156 => 
        N_156, N_1451_i => N_1451_i, N_1447_i => N_1447_i, 
        N_1452_i => N_1452_i, N_1446_i => N_1446_i, 
        wready_m_xhdl2 => wready_m_xhdl2, N_73_i_0 => N_73_i_0, 
        N_72_i => N_72_i, N_1445_i => N_1445_i, N_48 => N_48, 
        N_75_i => N_75_i, ahb_wr_done_sync => ahb_wr_done_sync, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, N_98 => N_98, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, araddr_arvalid_clr_d
         => araddr_arvalid_clr_d, awaddr_awvalid_clr_d => 
        awaddr_awvalid_clr_d, ahb_rd_req_sync => ahb_rd_req_sync, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID, latch_ahb_sig_sync
         => latch_ahb_sig_sync, 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, rdch_fifo_wr_en_r => 
        rdch_fifo_wr_en_r, COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, axi_read_rlast => 
        axi_read_rlast, HMASTLOCK_d => HMASTLOCK_d, HWRITE_d => 
        HWRITE_d, SDRCLK_c => SDRCLK_c, ARESET_n => ARESET_n);
    
    U_AHBAccCntrl : CoreAHBLtoAXI_AHBAccessControlHX
      port map(CoreAHBLite_0_AHBmslave10_HADDR(27) => 
        CoreAHBLite_0_AHBmslave10_HADDR(27), 
        CoreAHBLite_0_AHBmslave10_HADDR(26) => 
        CoreAHBLite_0_AHBmslave10_HADDR(26), 
        CoreAHBLite_0_AHBmslave10_HADDR(25) => 
        CoreAHBLite_0_AHBmslave10_HADDR(25), 
        CoreAHBLite_0_AHBmslave10_HADDR(24) => 
        CoreAHBLite_0_AHBmslave10_HADDR(24), 
        CoreAHBLite_0_AHBmslave10_HADDR(23) => 
        CoreAHBLite_0_AHBmslave10_HADDR(23), 
        CoreAHBLite_0_AHBmslave10_HADDR(22) => 
        CoreAHBLite_0_AHBmslave10_HADDR(22), 
        CoreAHBLite_0_AHBmslave10_HADDR(21) => 
        CoreAHBLite_0_AHBmslave10_HADDR(21), 
        CoreAHBLite_0_AHBmslave10_HADDR(20) => 
        CoreAHBLite_0_AHBmslave10_HADDR(20), 
        CoreAHBLite_0_AHBmslave10_HADDR(19) => 
        CoreAHBLite_0_AHBmslave10_HADDR(19), 
        CoreAHBLite_0_AHBmslave10_HADDR(18) => 
        CoreAHBLite_0_AHBmslave10_HADDR(18), 
        CoreAHBLite_0_AHBmslave10_HADDR(17) => 
        CoreAHBLite_0_AHBmslave10_HADDR(17), 
        CoreAHBLite_0_AHBmslave10_HADDR(16) => 
        CoreAHBLite_0_AHBmslave10_HADDR(16), 
        CoreAHBLite_0_AHBmslave10_HADDR(15) => 
        CoreAHBLite_0_AHBmslave10_HADDR(15), 
        CoreAHBLite_0_AHBmslave10_HADDR(14) => 
        CoreAHBLite_0_AHBmslave10_HADDR(14), 
        CoreAHBLite_0_AHBmslave10_HADDR(13) => 
        CoreAHBLite_0_AHBmslave10_HADDR(13), 
        CoreAHBLite_0_AHBmslave10_HADDR(12) => 
        CoreAHBLite_0_AHBmslave10_HADDR(12), 
        CoreAHBLite_0_AHBmslave10_HADDR(11) => 
        CoreAHBLite_0_AHBmslave10_HADDR(11), 
        CoreAHBLite_0_AHBmslave10_HADDR(10) => 
        CoreAHBLite_0_AHBmslave10_HADDR(10), 
        CoreAHBLite_0_AHBmslave10_HADDR(9) => 
        CoreAHBLite_0_AHBmslave10_HADDR(9), 
        CoreAHBLite_0_AHBmslave10_HADDR(8) => 
        CoreAHBLite_0_AHBmslave10_HADDR(8), 
        CoreAHBLite_0_AHBmslave10_HADDR(7) => 
        CoreAHBLite_0_AHBmslave10_HADDR(7), 
        CoreAHBLite_0_AHBmslave10_HADDR(6) => 
        CoreAHBLite_0_AHBmslave10_HADDR(6), 
        CoreAHBLite_0_AHBmslave10_HADDR(5) => 
        CoreAHBLite_0_AHBmslave10_HADDR(5), 
        CoreAHBLite_0_AHBmslave10_HADDR(4) => 
        CoreAHBLite_0_AHBmslave10_HADDR(4), 
        CoreAHBLite_0_AHBmslave10_HADDR(3) => 
        CoreAHBLite_0_AHBmslave10_HADDR(3), 
        CoreAHBLite_0_AHBmslave10_HADDR(2) => 
        CoreAHBLite_0_AHBmslave10_HADDR(2), 
        CoreAHBLite_0_AHBmslave10_HADDR(1) => 
        CoreAHBLite_0_AHBmslave10_HADDR(1), 
        CoreAHBLite_0_AHBmslave10_HADDR(0) => 
        CoreAHBLite_0_AHBmslave10_HADDR(0), HADDR_d(27) => 
        \HADDR_d[27]\, HADDR_d(26) => \HADDR_d[26]\, HADDR_d(25)
         => \HADDR_d[25]\, HADDR_d(24) => \HADDR_d[24]\, 
        HADDR_d(23) => \HADDR_d[23]\, HADDR_d(22) => 
        \HADDR_d[22]\, HADDR_d(21) => \HADDR_d[21]\, HADDR_d(20)
         => \HADDR_d[20]\, HADDR_d(19) => \HADDR_d[19]\, 
        HADDR_d(18) => \HADDR_d[18]\, HADDR_d(17) => 
        \HADDR_d[17]\, HADDR_d(16) => \HADDR_d[16]\, HADDR_d(15)
         => \HADDR_d[15]\, HADDR_d(14) => \HADDR_d[14]\, 
        HADDR_d(13) => \HADDR_d[13]\, HADDR_d(12) => 
        \HADDR_d[12]\, HADDR_d(11) => \HADDR_d[11]\, HADDR_d(10)
         => \HADDR_d[10]\, HADDR_d(9) => \HADDR_d[9]\, HADDR_d(8)
         => \HADDR_d[8]\, HADDR_d(7) => \HADDR_d[7]\, HADDR_d(6)
         => \HADDR_d[6]\, HADDR_d(5) => \HADDR_d[5]\, HADDR_d(4)
         => \HADDR_d[4]\, HADDR_d(3) => \HADDR_d[3]\, HADDR_d(2)
         => \HADDR_d[2]\, HADDR_d(1) => \HADDR_d[1]\, HADDR_d(0)
         => \HADDR_d[0]\, CoreAHBLite_0_AHBmslave10_HSIZE(1) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(1), 
        CoreAHBLite_0_AHBmslave10_HSIZE(0) => 
        CoreAHBLite_0_AHBmslave10_HSIZE(0), HSIZE_d(1) => 
        \HSIZE_d[1]\, HSIZE_d(0) => \HSIZE_d[0]\, 
        rdch_read_data(31) => \rdch_read_data[31]\, 
        rdch_read_data(30) => \rdch_read_data[30]\, 
        rdch_read_data(29) => \rdch_read_data[29]\, 
        rdch_read_data(28) => \rdch_read_data[28]\, 
        rdch_read_data(27) => \rdch_read_data[27]\, 
        rdch_read_data(26) => \rdch_read_data[26]\, 
        rdch_read_data(25) => \rdch_read_data[25]\, 
        rdch_read_data(24) => \rdch_read_data[24]\, 
        rdch_read_data(23) => \rdch_read_data[23]\, 
        rdch_read_data(22) => \rdch_read_data[22]\, 
        rdch_read_data(21) => \rdch_read_data[21]\, 
        rdch_read_data(20) => \rdch_read_data[20]\, 
        rdch_read_data(19) => \rdch_read_data[19]\, 
        rdch_read_data(18) => \rdch_read_data[18]\, 
        rdch_read_data(17) => \rdch_read_data[17]\, 
        rdch_read_data(16) => \rdch_read_data[16]\, 
        rdch_read_data(15) => \rdch_read_data[15]\, 
        rdch_read_data(14) => \rdch_read_data[14]\, 
        rdch_read_data(13) => \rdch_read_data[13]\, 
        rdch_read_data(12) => \rdch_read_data[12]\, 
        rdch_read_data(11) => \rdch_read_data[11]\, 
        rdch_read_data(10) => \rdch_read_data[10]\, 
        rdch_read_data(9) => \rdch_read_data[9]\, 
        rdch_read_data(8) => \rdch_read_data[8]\, 
        rdch_read_data(7) => \rdch_read_data[7]\, 
        rdch_read_data(6) => \rdch_read_data[6]\, 
        rdch_read_data(5) => \rdch_read_data[5]\, 
        rdch_read_data(4) => \rdch_read_data[4]\, 
        rdch_read_data(3) => \rdch_read_data[3]\, 
        rdch_read_data(2) => \rdch_read_data[2]\, 
        rdch_read_data(1) => \rdch_read_data[1]\, 
        rdch_read_data(0) => \rdch_read_data[0]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(31) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(31), 
        CoreAHBLite_0_AHBmslave10_HRDATA(30) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(30), 
        CoreAHBLite_0_AHBmslave10_HRDATA(29) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(29), 
        CoreAHBLite_0_AHBmslave10_HRDATA(28) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(28), 
        CoreAHBLite_0_AHBmslave10_HRDATA(27) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(27), 
        CoreAHBLite_0_AHBmslave10_HRDATA(26) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(26), 
        CoreAHBLite_0_AHBmslave10_HRDATA(25) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(25), 
        CoreAHBLite_0_AHBmslave10_HRDATA(24) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(24), 
        CoreAHBLite_0_AHBmslave10_HRDATA(23) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(23), 
        CoreAHBLite_0_AHBmslave10_HRDATA(22) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(22), 
        CoreAHBLite_0_AHBmslave10_HRDATA(21) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(21), 
        CoreAHBLite_0_AHBmslave10_HRDATA(20) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(20), 
        CoreAHBLite_0_AHBmslave10_HRDATA(19) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(19), 
        CoreAHBLite_0_AHBmslave10_HRDATA(18) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(18), 
        CoreAHBLite_0_AHBmslave10_HRDATA(17) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(17), 
        CoreAHBLite_0_AHBmslave10_HRDATA(16) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(16), 
        CoreAHBLite_0_AHBmslave10_HRDATA(15) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(15), 
        CoreAHBLite_0_AHBmslave10_HRDATA(14) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(14), 
        CoreAHBLite_0_AHBmslave10_HRDATA(13) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(13), 
        CoreAHBLite_0_AHBmslave10_HRDATA(12) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(12), 
        CoreAHBLite_0_AHBmslave10_HRDATA(11) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(11), 
        CoreAHBLite_0_AHBmslave10_HRDATA(10) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(10), 
        CoreAHBLite_0_AHBmslave10_HRDATA(9) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(9), 
        CoreAHBLite_0_AHBmslave10_HRDATA(8) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(8), 
        CoreAHBLite_0_AHBmslave10_HRDATA(7) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(7), 
        CoreAHBLite_0_AHBmslave10_HRDATA(6) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(6), 
        CoreAHBLite_0_AHBmslave10_HRDATA(5) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(5), 
        CoreAHBLite_0_AHBmslave10_HRDATA(4) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(4), 
        CoreAHBLite_0_AHBmslave10_HRDATA(3) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(3), 
        CoreAHBLite_0_AHBmslave10_HRDATA(2) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(2), 
        CoreAHBLite_0_AHBmslave10_HRDATA(1) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(1), 
        CoreAHBLite_0_AHBmslave10_HRDATA(0) => 
        CoreAHBLite_0_AHBmslave10_HRDATA(0), 
        CoreAHBLite_0_AHBmslave10_HWDATA(31) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(31), 
        CoreAHBLite_0_AHBmslave10_HWDATA(30) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(30), 
        CoreAHBLite_0_AHBmslave10_HWDATA(29) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(29), 
        CoreAHBLite_0_AHBmslave10_HWDATA(28) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(28), 
        CoreAHBLite_0_AHBmslave10_HWDATA(27) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(27), 
        CoreAHBLite_0_AHBmslave10_HWDATA(26) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(26), 
        CoreAHBLite_0_AHBmslave10_HWDATA(25) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(25), 
        CoreAHBLite_0_AHBmslave10_HWDATA(24) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(24), 
        CoreAHBLite_0_AHBmslave10_HWDATA(23) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(23), 
        CoreAHBLite_0_AHBmslave10_HWDATA(22) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(22), 
        CoreAHBLite_0_AHBmslave10_HWDATA(21) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(21), 
        CoreAHBLite_0_AHBmslave10_HWDATA(20) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(20), 
        CoreAHBLite_0_AHBmslave10_HWDATA(19) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(19), 
        CoreAHBLite_0_AHBmslave10_HWDATA(18) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(18), 
        CoreAHBLite_0_AHBmslave10_HWDATA(17) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(17), 
        CoreAHBLite_0_AHBmslave10_HWDATA(16) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(16), 
        CoreAHBLite_0_AHBmslave10_HWDATA(15) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(15), 
        CoreAHBLite_0_AHBmslave10_HWDATA(14) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(14), 
        CoreAHBLite_0_AHBmslave10_HWDATA(13) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(13), 
        CoreAHBLite_0_AHBmslave10_HWDATA(12) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(12), 
        CoreAHBLite_0_AHBmslave10_HWDATA(11) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(11), 
        CoreAHBLite_0_AHBmslave10_HWDATA(10) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(10), 
        CoreAHBLite_0_AHBmslave10_HWDATA(9) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(9), 
        CoreAHBLite_0_AHBmslave10_HWDATA(8) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(8), 
        CoreAHBLite_0_AHBmslave10_HWDATA(7) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(7), 
        CoreAHBLite_0_AHBmslave10_HWDATA(6) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(6), 
        CoreAHBLite_0_AHBmslave10_HWDATA(5) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(5), 
        CoreAHBLite_0_AHBmslave10_HWDATA(4) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(4), 
        CoreAHBLite_0_AHBmslave10_HWDATA(3) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(3), 
        CoreAHBLite_0_AHBmslave10_HWDATA(2) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(2), 
        CoreAHBLite_0_AHBmslave10_HWDATA(1) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(1), 
        CoreAHBLite_0_AHBmslave10_HWDATA(0) => 
        CoreAHBLite_0_AHBmslave10_HWDATA(0), wrch_hwdata_r(31)
         => \wrch_hwdata_r[31]\, wrch_hwdata_r(30) => 
        \wrch_hwdata_r[30]\, wrch_hwdata_r(29) => 
        \wrch_hwdata_r[29]\, wrch_hwdata_r(28) => 
        \wrch_hwdata_r[28]\, wrch_hwdata_r(27) => 
        \wrch_hwdata_r[27]\, wrch_hwdata_r(26) => 
        \wrch_hwdata_r[26]\, wrch_hwdata_r(25) => 
        \wrch_hwdata_r[25]\, wrch_hwdata_r(24) => 
        \wrch_hwdata_r[24]\, wrch_hwdata_r(23) => 
        \wrch_hwdata_r[23]\, wrch_hwdata_r(22) => 
        \wrch_hwdata_r[22]\, wrch_hwdata_r(21) => 
        \wrch_hwdata_r[21]\, wrch_hwdata_r(20) => 
        \wrch_hwdata_r[20]\, wrch_hwdata_r(19) => 
        \wrch_hwdata_r[19]\, wrch_hwdata_r(18) => 
        \wrch_hwdata_r[18]\, wrch_hwdata_r(17) => 
        \wrch_hwdata_r[17]\, wrch_hwdata_r(16) => 
        \wrch_hwdata_r[16]\, wrch_hwdata_r(15) => 
        \wrch_hwdata_r[15]\, wrch_hwdata_r(14) => 
        \wrch_hwdata_r[14]\, wrch_hwdata_r(13) => 
        \wrch_hwdata_r[13]\, wrch_hwdata_r(12) => 
        \wrch_hwdata_r[12]\, wrch_hwdata_r(11) => 
        \wrch_hwdata_r[11]\, wrch_hwdata_r(10) => 
        \wrch_hwdata_r[10]\, wrch_hwdata_r(9) => 
        \wrch_hwdata_r[9]\, wrch_hwdata_r(8) => 
        \wrch_hwdata_r[8]\, wrch_hwdata_r(7) => 
        \wrch_hwdata_r[7]\, wrch_hwdata_r(6) => 
        \wrch_hwdata_r[6]\, wrch_hwdata_r(5) => 
        \wrch_hwdata_r[5]\, wrch_hwdata_r(4) => 
        \wrch_hwdata_r[4]\, wrch_hwdata_r(3) => 
        \wrch_hwdata_r[3]\, wrch_hwdata_r(2) => 
        \wrch_hwdata_r[2]\, wrch_hwdata_r(1) => 
        \wrch_hwdata_r[1]\, wrch_hwdata_r(0) => 
        \wrch_hwdata_r[0]\, xhdl1222_0 => xhdl1222_0, 
        synchronizer_1_0 => \synchronizer_1[0]\, 
        masterAddrInProg_0 => masterAddrInProg_0, current_state_0
         => current_state_0, N_92 => N_92, m0PrevDataSlaveReady
         => m0PrevDataSlaveReady, N_91 => N_91, post_sync_1_reg
         => post_sync_1_reg, rdch_fifo_empty => rdch_fifo_empty, 
        N_163_i => N_163_i, hsel2 => hsel2, hsel2_0_a2_1 => 
        hsel2_0_a2_1, valid_ahbcmd_i_o3_1 => valid_ahbcmd_i_o3_1, 
        rdch_fifo_rd_en_r => rdch_fifo_rd_en_r, latch_ahb_sig => 
        latch_ahb_sig, BVALID_sync => BVALID_sync, ahb_wr_done
         => ahb_wr_done, CoreAHBLite_0_AHBmslave10_HMASTLOCK => 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, HMASTLOCK_d => 
        HMASTLOCK_d, CoreAHBLite_0_AHBmslave10_HWRITE => 
        CoreAHBLite_0_AHBmslave10_HWRITE, HWRITE_d => HWRITE_d, 
        SDRCLK_c => SDRCLK_c, ARESET_n => ARESET_n, 
        ahb_busyidle_cyc_i => ahb_busyidle_cyc_i, 
        ahb_busyidle_cyc => ahb_busyidle_cyc);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top_sb is

    port( DQ_in              : in    std_logic_vector(15 downto 0);
          BA_c               : out   std_logic_vector(1 downto 0);
          SA_c               : out   std_logic_vector(11 downto 0);
          sdr_datain_reg     : out   std_logic_vector(15 downto 0);
          DQM_c              : out   std_logic_vector(1 downto 0);
          CS_N_c_0           : out   std_logic;
          CAS_N_c            : out   std_logic;
          CKE_c              : out   std_logic;
          un1_top_sb_0_3_i_i : out   std_logic;
          RAS_N_c            : out   std_logic;
          WE_N_c             : out   std_logic;
          SPI_0_SS0          : inout std_logic := 'Z';
          SPI_0_DO           : out   std_logic;
          SPI_0_DI           : in    std_logic;
          SPI_0_CLK          : inout std_logic := 'Z';
          MMUART_0_TXD       : out   std_logic;
          MMUART_0_RXD       : in    std_logic;
          I2C_0_SDA          : inout std_logic := 'Z';
          I2C_0_SCL          : inout std_logic := 'Z';
          GPIO_29_BI         : inout std_logic := 'Z';
          GPIO_26_BI         : inout std_logic := 'Z';
          GPIO_25_BI         : inout std_logic := 'Z';
          GPIO_24_BI         : inout std_logic := 'Z';
          GPIO_23_BI         : inout std_logic := 'Z';
          GPIO_22_BI         : inout std_logic := 'Z';
          GPIO_21_BI         : inout std_logic := 'Z';
          GPIO_20_BI         : inout std_logic := 'Z';
          GPIO_19_BI         : inout std_logic := 'Z';
          GPIO_18_BI         : inout std_logic := 'Z';
          GPIO_17_BI         : inout std_logic := 'Z';
          GPIO_16_BI         : inout std_logic := 'Z';
          GPIO_15_BI         : inout std_logic := 'Z';
          GPIO_14_BI         : inout std_logic := 'Z';
          GPIO_13_BI         : inout std_logic := 'Z';
          GPIO_12_BI         : inout std_logic := 'Z';
          GPIO_11_BI         : inout std_logic := 'Z';
          GPIO_10_BI         : inout std_logic := 'Z';
          GPIO_9_BI          : inout std_logic := 'Z';
          GPIO_8_BI          : inout std_logic := 'Z';
          GPIO_1_BI          : inout std_logic := 'Z';
          CAN_TX             : out   std_logic;
          CAN_TX_EN_N        : out   std_logic;
          CAN_RX             : in    std_logic;
          SDRCLK_c           : out   std_logic;
          CLK1_PAD           : in    std_logic;
          DEVRST_N           : in    std_logic
        );

end top_sb;

architecture DEF_ARCH of top_sb is 

  component CORESDR_AXI
    port( COREAXI_0_AXImslave16_AWSIZE       : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_ARSIZE       : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_WDATA        : in    std_logic_vector(63 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_AWADDR       : in    std_logic_vector(23 downto 1) := (others => 'U');
          COREAXI_0_AXImslave16_ARADDR       : in    std_logic_vector(23 downto 1) := (others => 'U');
          COREAXI_0_AXImslave16_WSTRB        : in    std_logic_vector(7 downto 0) := (others => 'U');
          DQM_c                              : out   std_logic_vector(1 downto 0);
          sdr_datain_reg                     : out   std_logic_vector(15 downto 0);
          SA_c                               : out   std_logic_vector(11 downto 0);
          BA_c                               : out   std_logic_vector(1 downto 0);
          DQ_in                              : in    std_logic_vector(15 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_RDATA_m_8    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_11   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_12   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_13   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_14   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_15   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_0    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_4    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_5    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_6    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_7    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_10   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_9    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_1    : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_34   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_47   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_19   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_20   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_21   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_23   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_41   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_33   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_42   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_49   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_50   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_57   : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_m_58   : out   std_logic;
          COREAXI_0_AXImslave16_ARBURST_0    : in    std_logic := 'U';
          CS_N_c_0                           : out   std_logic;
          axi_state_0                        : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_0      : out   std_logic;
          COREAXI_0_AXImslave16_RDATA_3      : out   std_logic;
          RDATA_reg_0                        : out   std_logic;
          RDATA_reg_3                        : out   std_logic;
          N_8_i                              : out   std_logic;
          N_23                               : in    std_logic := 'U';
          N_3169_i                           : out   std_logic;
          N_77_mux_i                         : out   std_logic;
          N_76_mux_i                         : out   std_logic;
          N_75_mux_i                         : out   std_logic;
          N_69_mux_i                         : out   std_logic;
          N_68_mux_i                         : out   std_logic;
          N_67_mux_i                         : out   std_logic;
          N_72_mux_i                         : out   std_logic;
          N_71_mux_i                         : out   std_logic;
          N_70_mux_i                         : out   std_logic;
          N_80_mux_i                         : out   std_logic;
          N_79_mux_i                         : out   std_logic;
          N_78_mux_i                         : out   std_logic;
          N_3297                             : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID : in    std_logic := 'U';
          N_3170_i                           : out   std_logic;
          COREAXI_0_AXImslave16_AWVALID      : in    std_logic := 'U';
          N_39                               : out   std_logic;
          WREADY_SI16_i                      : out   std_logic;
          COREAXI_0_AXImslave16_WVALID       : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID      : in    std_logic := 'U';
          i22_mux_2_i                        : out   std_logic;
          i22_mux_3_i                        : out   std_logic;
          i22_mux_4_i                        : out   std_logic;
          i22_mux_5_i                        : out   std_logic;
          i17_mux_2_i                        : out   std_logic;
          i17_mux_i                          : out   std_logic;
          i17_mux_0_i                        : out   std_logic;
          i17_mux_1_i                        : out   std_logic;
          i22_mux_i                          : out   std_logic;
          i22_mux_0_i                        : out   std_logic;
          i22_mux_1_i                        : out   std_logic;
          N_389                              : out   std_logic;
          N_3064_i                           : out   std_logic;
          N_3066_i                           : out   std_logic;
          N_3092_i                           : out   std_logic;
          N_3094_i                           : out   std_logic;
          N_3096_i                           : out   std_logic;
          N_3098_i                           : out   std_logic;
          N_3100_i                           : out   std_logic;
          N_3102_i                           : out   std_logic;
          N_74                               : out   std_logic;
          N_3167_i                           : in    std_logic := 'U';
          WE_N_c                             : out   std_logic;
          RAS_N_c                            : out   std_logic;
          un1_top_sb_0_3_i_i                 : out   std_logic;
          CKE_c                              : out   std_logic;
          CAS_N_c                            : out   std_logic;
          COREAXI_0_AXImslave16_BVALID       : out   std_logic;
          COREAXI_0_AXImslave16_AWREADY      : out   std_logic;
          COREAXI_0_AXImslave16_ARREADY      : out   std_logic;
          WREADY_SI16                        : out   std_logic;
          SDRCLK_c                           : in    std_logic := 'U';
          MSS_READY                          : in    std_logic := 'U'
        );
  end component;

  component CoreResetP
    port( top_sb_0_POWER_ON_RESET_N             : in    std_logic := 'U';
          top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MSS_RESET_N_M2F      : in    std_logic := 'U';
          CORERESETP_0_RESET_N_F2M              : out   std_logic;
          SDRCLK_c                              : in    std_logic := 'U';
          MSS_READY                             : out   std_logic
        );
  end component;

  component CoreAHBLite
    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : in    std_logic_vector(31 downto 0) := (others => 'U');
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HADDR               : out   std_logic_vector(27 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE               : out   std_logic_vector(1 downto 0);
          CoreAHBLite_0_AHBmslave10_HWDATA              : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : in    std_logic_vector(31 downto 0) := (others => 'U');
          masterAddrInProg_0                            : out   std_logic;
          current_state_0                               : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : out   std_logic;
          xhdl1222_0                                    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : out   std_logic;
          N_92                                          : out   std_logic;
          N_91                                          : out   std_logic;
          hready_m_xhdl349                              : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : in    std_logic := 'U';
          m0PrevDataSlaveReady                          : out   std_logic;
          SDRCLK_c                                      : in    std_logic := 'U';
          MSS_READY                                     : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave10_HMASTLOCK           : out   std_logic;
          CoreAHBLite_0_AHBmslave10_HWRITE              : out   std_logic;
          hsel2                                         : out   std_logic;
          hsel2_0_a2_1                                  : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component top_sb_CCC_0_FCCC
    port( FAB_CCC_LOCK : out   std_logic;
          CLK1_PAD     : in    std_logic := 'U';
          SDRCLK_c     : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component top_sb_MSS
    port( top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE    : out   std_logic_vector(1 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA   : out   std_logic_vector(31 downto 0);
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR    : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HRDATA              : in    std_logic_vector(31 downto 0) := (others => 'U');
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0  : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY   : in    std_logic := 'U';
          SDRCLK_c                                      : in    std_logic := 'U';
          CORERESETP_0_RESET_N_F2M                      : in    std_logic := 'U';
          FAB_CCC_LOCK                                  : in    std_logic := 'U';
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK    : out   std_logic;
          top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE   : out   std_logic;
          top_sb_MSS_TMP_0_MSS_RESET_N_M2F              : out   std_logic;
          top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N         : out   std_logic;
          hready_m_xhdl349                              : in    std_logic := 'U';
          CAN_RX                                        : in    std_logic := 'U';
          CAN_TX_EN_N                                   : out   std_logic;
          CAN_TX                                        : out   std_logic;
          GPIO_1_BI                                     : inout   std_logic;
          GPIO_8_BI                                     : inout   std_logic;
          GPIO_9_BI                                     : inout   std_logic;
          GPIO_10_BI                                    : inout   std_logic;
          GPIO_11_BI                                    : inout   std_logic;
          GPIO_12_BI                                    : inout   std_logic;
          GPIO_13_BI                                    : inout   std_logic;
          GPIO_14_BI                                    : inout   std_logic;
          GPIO_15_BI                                    : inout   std_logic;
          GPIO_16_BI                                    : inout   std_logic;
          GPIO_17_BI                                    : inout   std_logic;
          GPIO_18_BI                                    : inout   std_logic;
          GPIO_19_BI                                    : inout   std_logic;
          GPIO_20_BI                                    : inout   std_logic;
          GPIO_21_BI                                    : inout   std_logic;
          GPIO_22_BI                                    : inout   std_logic;
          GPIO_23_BI                                    : inout   std_logic;
          GPIO_24_BI                                    : inout   std_logic;
          GPIO_25_BI                                    : inout   std_logic;
          GPIO_26_BI                                    : inout   std_logic;
          GPIO_29_BI                                    : inout   std_logic;
          I2C_0_SCL                                     : inout   std_logic;
          I2C_0_SDA                                     : inout   std_logic;
          MMUART_0_RXD                                  : in    std_logic := 'U';
          MMUART_0_TXD                                  : out   std_logic;
          SPI_0_CLK                                     : inout   std_logic;
          SPI_0_DI                                      : in    std_logic := 'U';
          SPI_0_DO                                      : out   std_logic;
          SPI_0_SS0                                     : inout   std_logic
        );
  end component;

  component top_sb_COREAXI_0_COREAXI
    port( COREAXI_0_AXImslave16_AWSIZE         : out   std_logic_vector(1 downto 0);
          COREAXI_0_AXImslave16_ARADDR         : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_AWADDR         : out   std_logic_vector(23 downto 1);
          COREAXI_0_AXImslave16_WSTRB          : out   std_logic_vector(7 downto 0);
          COREAXI_0_AXImslave16_WDATA          : out   std_logic_vector(63 downto 0);
          COREAXI_0_AXImslave16_ARSIZE         : out   std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : out   std_logic_vector(63 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : in    std_logic_vector(63 downto 16) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : in    std_logic_vector(27 downto 1) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : in    std_logic_vector(1 downto 0) := (others => 'U');
          COREAXI_0_AXImslave16_ARBURST_0      : out   std_logic;
          axi_current_state_0                  : in    std_logic := 'U';
          axi_current_state_3                  : in    std_logic := 'U';
          axi_state_0                          : in    std_logic := 'U';
          RDATA_reg_3                          : in    std_logic := 'U';
          RDATA_reg_0                          : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_3        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_0        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_57     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_58     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_41     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_42     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_47     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_49     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_50     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_33     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_34     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_11     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_12     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_13     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_14     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_15     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_19     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_20     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_21     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_23     : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_0      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_1      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_4      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_5      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_6      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_7      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_8      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_9      : in    std_logic := 'U';
          COREAXI_0_AXImslave16_RDATA_m_10     : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : in    std_logic := 'U';
          COREAXI_0_AXImslave16_WVALID         : out   std_logic;
          WREADY_SI16_i                        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_AWVALID        : out   std_logic;
          COREAXI_0_AXImslave16_AWREADY        : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : out   std_logic;
          wready_m_xhdl2                       : out   std_logic;
          N_1445_i                             : in    std_logic := 'U';
          N_1446_i                             : in    std_logic := 'U';
          N_1447_i                             : in    std_logic := 'U';
          N_1448_i                             : in    std_logic := 'U';
          N_1449_i                             : in    std_logic := 'U';
          N_1450_i                             : in    std_logic := 'U';
          N_1451_i                             : in    std_logic := 'U';
          N_1452_i                             : in    std_logic := 'U';
          N_202_i                              : in    std_logic := 'U';
          N_201_i                              : in    std_logic := 'U';
          N_200_i                              : in    std_logic := 'U';
          N_197_i                              : in    std_logic := 'U';
          N_195_i                              : in    std_logic := 'U';
          N_134_i                              : in    std_logic := 'U';
          N_133_i                              : in    std_logic := 'U';
          N_380_i                              : in    std_logic := 'U';
          N_278_i                              : in    std_logic := 'U';
          N_381_i                              : in    std_logic := 'U';
          N_382_i                              : in    std_logic := 'U';
          N_277_i                              : in    std_logic := 'U';
          N_276_i                              : in    std_logic := 'U';
          N_275_i                              : in    std_logic := 'U';
          N_274_i                              : in    std_logic := 'U';
          N_273_i                              : in    std_logic := 'U';
          N_272_i                              : in    std_logic := 'U';
          N_203_i                              : in    std_logic := 'U';
          N_137_i                              : in    std_logic := 'U';
          N_136_i                              : in    std_logic := 'U';
          N_135_i                              : in    std_logic := 'U';
          N_48                                 : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : out   std_logic;
          araddr_arvalid_clr_d                 : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : in    std_logic := 'U';
          awaddr_awvalid_clr_d                 : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          COREAXI_0_AXImslave16_BVALID         : in    std_logic := 'U';
          N_3297                               : in    std_logic := 'U';
          N_389                                : in    std_logic := 'U';
          N_74                                 : in    std_logic := 'U';
          N_3167_i                             : out   std_logic;
          N_23                                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : in    std_logic := 'U';
          N_3170_i                             : in    std_logic := 'U';
          N_39                                 : in    std_logic := 'U';
          N_78_mux_i                           : in    std_logic := 'U';
          N_79_mux_i                           : in    std_logic := 'U';
          N_80_mux_i                           : in    std_logic := 'U';
          N_70_mux_i                           : in    std_logic := 'U';
          N_71_mux_i                           : in    std_logic := 'U';
          N_72_mux_i                           : in    std_logic := 'U';
          N_3094_i                             : in    std_logic := 'U';
          N_3096_i                             : in    std_logic := 'U';
          N_3098_i                             : in    std_logic := 'U';
          N_3100_i                             : in    std_logic := 'U';
          N_3102_i                             : in    std_logic := 'U';
          N_3169_i                             : in    std_logic := 'U';
          N_3066_i                             : in    std_logic := 'U';
          N_67_mux_i                           : in    std_logic := 'U';
          N_68_mux_i                           : in    std_logic := 'U';
          N_69_mux_i                           : in    std_logic := 'U';
          N_75_mux_i                           : in    std_logic := 'U';
          N_76_mux_i                           : in    std_logic := 'U';
          N_77_mux_i                           : in    std_logic := 'U';
          i22_mux_2_i                          : in    std_logic := 'U';
          i22_mux_3_i                          : in    std_logic := 'U';
          i22_mux_4_i                          : in    std_logic := 'U';
          i22_mux_5_i                          : in    std_logic := 'U';
          N_8_i                                : in    std_logic := 'U';
          i17_mux_2_i                          : in    std_logic := 'U';
          N_3064_i                             : in    std_logic := 'U';
          N_3092_i                             : in    std_logic := 'U';
          i17_mux_i                            : in    std_logic := 'U';
          i17_mux_0_i                          : in    std_logic := 'U';
          i17_mux_1_i                          : in    std_logic := 'U';
          i22_mux_i                            : in    std_logic := 'U';
          i22_mux_0_i                          : in    std_logic := 'U';
          i22_mux_1_i                          : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARREADY        : in    std_logic := 'U';
          COREAXI_0_AXImslave16_ARVALID        : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : in    std_logic := 'U';
          WREADY_SI16                          : in    std_logic := 'U';
          N_75_i                               : in    std_logic := 'U'
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI
    port( COREAHBLTOAXI_0_AXIMasterIF_ARSIZE   : out   std_logic_vector(1 downto 0);
          COREAHBLTOAXI_0_AXIMasterIF_ARADDR   : out   std_logic_vector(27 downto 1);
          COREAHBLTOAXI_0_AXIMasterIF_RDATA    : in    std_logic_vector(63 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_WDATA    : out   std_logic_vector(63 downto 16);
          CoreAHBLite_0_AHBmslave10_HWDATA     : in    std_logic_vector(31 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HRDATA     : out   std_logic_vector(31 downto 0);
          CoreAHBLite_0_AHBmslave10_HSIZE      : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAHBLite_0_AHBmslave10_HADDR      : in    std_logic_vector(27 downto 0) := (others => 'U');
          COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 : out   std_logic;
          axi_current_state_0                  : out   std_logic;
          axi_current_state_3                  : out   std_logic;
          current_state_0                      : out   std_logic;
          masterAddrInProg_0                   : in    std_logic := 'U';
          xhdl1222_0                           : in    std_logic := 'U';
          MSS_READY                            : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RREADY   : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WVALID   : out   std_logic;
          awaddr_awvalid_clr_d                 : out   std_logic;
          araddr_arvalid_clr_d                 : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_WREADY   : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_AWREADY  : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RVALID   : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_RLAST    : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARREADY  : in    std_logic := 'U';
          COREAHBLTOAXI_0_AXIMasterIF_ARVALID  : out   std_logic;
          N_75_i                               : out   std_logic;
          N_48                                 : out   std_logic;
          N_1445_i                             : out   std_logic;
          wready_m_xhdl2                       : in    std_logic := 'U';
          N_1446_i                             : out   std_logic;
          N_1452_i                             : out   std_logic;
          N_1447_i                             : out   std_logic;
          N_1451_i                             : out   std_logic;
          N_135_i                              : out   std_logic;
          N_136_i                              : out   std_logic;
          N_137_i                              : out   std_logic;
          N_203_i                              : out   std_logic;
          N_272_i                              : out   std_logic;
          N_273_i                              : out   std_logic;
          N_274_i                              : out   std_logic;
          N_275_i                              : out   std_logic;
          N_276_i                              : out   std_logic;
          N_277_i                              : out   std_logic;
          N_382_i                              : out   std_logic;
          N_381_i                              : out   std_logic;
          N_278_i                              : out   std_logic;
          N_380_i                              : out   std_logic;
          N_133_i                              : out   std_logic;
          N_134_i                              : out   std_logic;
          N_195_i                              : out   std_logic;
          N_197_i                              : out   std_logic;
          N_200_i                              : out   std_logic;
          N_201_i                              : out   std_logic;
          N_202_i                              : out   std_logic;
          N_1450_i                             : out   std_logic;
          N_1449_i                             : out   std_logic;
          N_1448_i                             : out   std_logic;
          COREAHBLTOAXI_0_AXIMasterIF_BVALID   : in    std_logic := 'U';
          SDRCLK_c                             : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave10_HWRITE     : in    std_logic := 'U';
          CoreAHBLite_0_AHBmslave10_HMASTLOCK  : in    std_logic := 'U';
          hsel2_0_a2_1                         : in    std_logic := 'U';
          hsel2                                : in    std_logic := 'U';
          N_91                                 : in    std_logic := 'U';
          m0PrevDataSlaveReady                 : in    std_logic := 'U';
          N_92                                 : in    std_logic := 'U'
        );
  end component;

    signal top_sb_0_POWER_ON_RESET_N, FAB_CCC_LOCK, \SDRCLK_c\, 
        \masterAddrInProg[0]\, \current_state[7]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS[1]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP[0]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[0]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[1]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[2]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[3]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[4]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[5]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[6]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[7]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[8]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[9]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[10]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[11]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[12]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[13]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[14]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[15]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[16]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[17]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[18]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[19]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[20]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[21]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[22]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[23]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[24]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[25]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[26]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[27]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[28]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[29]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[30]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[31]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[0]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[1]\, 
        \xhdl1222[10]\, \CoreAHBLite_0_AHBmslave10_HADDR[0]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[1]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[2]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[3]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[4]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[5]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[6]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[7]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[8]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[9]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[10]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[11]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[12]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[13]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[14]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[15]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[16]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[17]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[18]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[19]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[20]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[21]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[22]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[23]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[24]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[25]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[26]\, 
        \CoreAHBLite_0_AHBmslave10_HADDR[27]\, 
        \CoreAHBLite_0_AHBmslave10_HSIZE[0]\, 
        \CoreAHBLite_0_AHBmslave10_HSIZE[1]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[0]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[1]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[2]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[3]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[4]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[5]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[6]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[7]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[8]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[9]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[10]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[11]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[12]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[13]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[14]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[15]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[16]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[17]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[18]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[19]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[20]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[21]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[22]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[23]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[24]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[25]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[26]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[27]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[28]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[29]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[30]\, 
        \CoreAHBLite_0_AHBmslave10_HWDATA[31]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[0]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[1]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[2]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[3]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[4]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[5]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[6]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[7]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[8]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[9]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[10]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[11]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[12]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[13]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[14]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[15]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[16]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[17]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[18]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[19]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[20]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[21]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[22]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[23]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[24]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[25]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[26]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[27]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[28]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[29]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[30]\, 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[31]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY, N_92, N_91, 
        hready_m_xhdl349, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        m0PrevDataSlaveReady, MSS_READY, 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, 
        CoreAHBLite_0_AHBmslave10_HWRITE, hsel2, hsel2_0_a2_1, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[3]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[4]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[5]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[6]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[7]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[8]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[9]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[10]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[11]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[12]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[13]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[14]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[15]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[16]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[17]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[18]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[19]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[20]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[21]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[22]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[23]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[24]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[25]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[26]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[27]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[0]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[1]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[2]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[3]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[4]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[5]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[6]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[7]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[8]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[9]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[10]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[11]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[12]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[13]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[14]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[15]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[16]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[17]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[18]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[19]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[20]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[21]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[22]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[23]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[24]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[25]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[26]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[27]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[28]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[29]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[30]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[31]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[32]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[33]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[34]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[35]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[36]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[37]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[38]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[39]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[40]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[41]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[42]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[43]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[44]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[45]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[46]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[47]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[48]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[49]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[50]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[51]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[52]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[53]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[54]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[55]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[56]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[57]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[58]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[59]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[60]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[61]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[62]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[63]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_ARLOCK[1]\, 
        \axi_current_state[1]\, \axi_current_state[4]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[16]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[17]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[18]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[22]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[23]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[24]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[25]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[26]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[27]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[29]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[30]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[32]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[33]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[34]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[35]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[36]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[37]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[38]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[39]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[40]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[41]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[42]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[43]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[44]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[45]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[46]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[47]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[48]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[49]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[50]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[51]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[52]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[53]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[54]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[55]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[56]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[57]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[58]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[59]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[60]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[61]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[62]\, 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[63]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[0]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[1]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[2]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[3]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[4]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[5]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[6]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[7]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[8]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[9]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[10]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[11]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[12]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[13]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[14]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[15]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[16]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[17]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[18]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[19]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[20]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[21]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[22]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[23]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[24]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[25]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[26]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[27]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[28]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[29]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[30]\, 
        \CoreAHBLite_0_AHBmslave10_HRDATA[31]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, awaddr_awvalid_clr_d, 
        araddr_arvalid_clr_d, COREAHBLTOAXI_0_AXIMasterIF_WREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, N_75_i, N_48, 
        N_1445_i, wready_m_xhdl2, N_1446_i, N_1452_i, N_1447_i, 
        N_1451_i, N_135_i, N_136_i, N_137_i, N_203_i, N_272_i, 
        N_273_i, N_274_i, N_275_i, N_276_i, N_277_i, N_382_i, 
        N_381_i, N_278_i, N_380_i, N_133_i, N_134_i, N_195_i, 
        N_197_i, N_200_i, N_201_i, N_202_i, N_1450_i, N_1449_i, 
        N_1448_i, COREAHBLTOAXI_0_AXIMasterIF_BVALID, 
        \COREAXI_0_AXImslave16_AWSIZE[0]\, 
        \COREAXI_0_AXImslave16_AWSIZE[1]\, 
        \COREAXI_0_AXImslave16_ARADDR[1]\, 
        \COREAXI_0_AXImslave16_ARADDR[2]\, 
        \COREAXI_0_AXImslave16_ARADDR[3]\, 
        \COREAXI_0_AXImslave16_ARADDR[4]\, 
        \COREAXI_0_AXImslave16_ARADDR[5]\, 
        \COREAXI_0_AXImslave16_ARADDR[6]\, 
        \COREAXI_0_AXImslave16_ARADDR[7]\, 
        \COREAXI_0_AXImslave16_ARADDR[8]\, 
        \COREAXI_0_AXImslave16_ARADDR[9]\, 
        \COREAXI_0_AXImslave16_ARADDR[10]\, 
        \COREAXI_0_AXImslave16_ARADDR[11]\, 
        \COREAXI_0_AXImslave16_ARADDR[12]\, 
        \COREAXI_0_AXImslave16_ARADDR[13]\, 
        \COREAXI_0_AXImslave16_ARADDR[14]\, 
        \COREAXI_0_AXImslave16_ARADDR[15]\, 
        \COREAXI_0_AXImslave16_ARADDR[16]\, 
        \COREAXI_0_AXImslave16_ARADDR[17]\, 
        \COREAXI_0_AXImslave16_ARADDR[18]\, 
        \COREAXI_0_AXImslave16_ARADDR[19]\, 
        \COREAXI_0_AXImslave16_ARADDR[20]\, 
        \COREAXI_0_AXImslave16_ARADDR[21]\, 
        \COREAXI_0_AXImslave16_ARADDR[22]\, 
        \COREAXI_0_AXImslave16_ARADDR[23]\, 
        \COREAXI_0_AXImslave16_AWADDR[1]\, 
        \COREAXI_0_AXImslave16_AWADDR[2]\, 
        \COREAXI_0_AXImslave16_AWADDR[3]\, 
        \COREAXI_0_AXImslave16_AWADDR[4]\, 
        \COREAXI_0_AXImslave16_AWADDR[5]\, 
        \COREAXI_0_AXImslave16_AWADDR[6]\, 
        \COREAXI_0_AXImslave16_AWADDR[7]\, 
        \COREAXI_0_AXImslave16_AWADDR[8]\, 
        \COREAXI_0_AXImslave16_AWADDR[9]\, 
        \COREAXI_0_AXImslave16_AWADDR[10]\, 
        \COREAXI_0_AXImslave16_AWADDR[11]\, 
        \COREAXI_0_AXImslave16_AWADDR[12]\, 
        \COREAXI_0_AXImslave16_AWADDR[13]\, 
        \COREAXI_0_AXImslave16_AWADDR[14]\, 
        \COREAXI_0_AXImslave16_AWADDR[15]\, 
        \COREAXI_0_AXImslave16_AWADDR[16]\, 
        \COREAXI_0_AXImslave16_AWADDR[17]\, 
        \COREAXI_0_AXImslave16_AWADDR[18]\, 
        \COREAXI_0_AXImslave16_AWADDR[19]\, 
        \COREAXI_0_AXImslave16_AWADDR[20]\, 
        \COREAXI_0_AXImslave16_AWADDR[21]\, 
        \COREAXI_0_AXImslave16_AWADDR[22]\, 
        \COREAXI_0_AXImslave16_AWADDR[23]\, 
        \COREAXI_0_AXImslave16_WSTRB[0]\, 
        \COREAXI_0_AXImslave16_WSTRB[1]\, 
        \COREAXI_0_AXImslave16_WSTRB[2]\, 
        \COREAXI_0_AXImslave16_WSTRB[3]\, 
        \COREAXI_0_AXImslave16_WSTRB[4]\, 
        \COREAXI_0_AXImslave16_WSTRB[5]\, 
        \COREAXI_0_AXImslave16_WSTRB[6]\, 
        \COREAXI_0_AXImslave16_WSTRB[7]\, 
        \COREAXI_0_AXImslave16_WDATA[0]\, 
        \COREAXI_0_AXImslave16_WDATA[1]\, 
        \COREAXI_0_AXImslave16_WDATA[2]\, 
        \COREAXI_0_AXImslave16_WDATA[3]\, 
        \COREAXI_0_AXImslave16_WDATA[4]\, 
        \COREAXI_0_AXImslave16_WDATA[5]\, 
        \COREAXI_0_AXImslave16_WDATA[6]\, 
        \COREAXI_0_AXImslave16_WDATA[7]\, 
        \COREAXI_0_AXImslave16_WDATA[8]\, 
        \COREAXI_0_AXImslave16_WDATA[9]\, 
        \COREAXI_0_AXImslave16_WDATA[10]\, 
        \COREAXI_0_AXImslave16_WDATA[11]\, 
        \COREAXI_0_AXImslave16_WDATA[12]\, 
        \COREAXI_0_AXImslave16_WDATA[13]\, 
        \COREAXI_0_AXImslave16_WDATA[14]\, 
        \COREAXI_0_AXImslave16_WDATA[15]\, 
        \COREAXI_0_AXImslave16_WDATA[16]\, 
        \COREAXI_0_AXImslave16_WDATA[17]\, 
        \COREAXI_0_AXImslave16_WDATA[18]\, 
        \COREAXI_0_AXImslave16_WDATA[19]\, 
        \COREAXI_0_AXImslave16_WDATA[20]\, 
        \COREAXI_0_AXImslave16_WDATA[21]\, 
        \COREAXI_0_AXImslave16_WDATA[22]\, 
        \COREAXI_0_AXImslave16_WDATA[23]\, 
        \COREAXI_0_AXImslave16_WDATA[24]\, 
        \COREAXI_0_AXImslave16_WDATA[25]\, 
        \COREAXI_0_AXImslave16_WDATA[26]\, 
        \COREAXI_0_AXImslave16_WDATA[27]\, 
        \COREAXI_0_AXImslave16_WDATA[28]\, 
        \COREAXI_0_AXImslave16_WDATA[29]\, 
        \COREAXI_0_AXImslave16_WDATA[30]\, 
        \COREAXI_0_AXImslave16_WDATA[31]\, 
        \COREAXI_0_AXImslave16_WDATA[32]\, 
        \COREAXI_0_AXImslave16_WDATA[33]\, 
        \COREAXI_0_AXImslave16_WDATA[34]\, 
        \COREAXI_0_AXImslave16_WDATA[35]\, 
        \COREAXI_0_AXImslave16_WDATA[36]\, 
        \COREAXI_0_AXImslave16_WDATA[37]\, 
        \COREAXI_0_AXImslave16_WDATA[38]\, 
        \COREAXI_0_AXImslave16_WDATA[39]\, 
        \COREAXI_0_AXImslave16_WDATA[40]\, 
        \COREAXI_0_AXImslave16_WDATA[41]\, 
        \COREAXI_0_AXImslave16_WDATA[42]\, 
        \COREAXI_0_AXImslave16_WDATA[43]\, 
        \COREAXI_0_AXImslave16_WDATA[44]\, 
        \COREAXI_0_AXImslave16_WDATA[45]\, 
        \COREAXI_0_AXImslave16_WDATA[46]\, 
        \COREAXI_0_AXImslave16_WDATA[47]\, 
        \COREAXI_0_AXImslave16_WDATA[48]\, 
        \COREAXI_0_AXImslave16_WDATA[49]\, 
        \COREAXI_0_AXImslave16_WDATA[50]\, 
        \COREAXI_0_AXImslave16_WDATA[51]\, 
        \COREAXI_0_AXImslave16_WDATA[52]\, 
        \COREAXI_0_AXImslave16_WDATA[53]\, 
        \COREAXI_0_AXImslave16_WDATA[54]\, 
        \COREAXI_0_AXImslave16_WDATA[55]\, 
        \COREAXI_0_AXImslave16_WDATA[56]\, 
        \COREAXI_0_AXImslave16_WDATA[57]\, 
        \COREAXI_0_AXImslave16_WDATA[58]\, 
        \COREAXI_0_AXImslave16_WDATA[59]\, 
        \COREAXI_0_AXImslave16_WDATA[60]\, 
        \COREAXI_0_AXImslave16_WDATA[61]\, 
        \COREAXI_0_AXImslave16_WDATA[62]\, 
        \COREAXI_0_AXImslave16_WDATA[63]\, 
        \COREAXI_0_AXImslave16_ARSIZE[0]\, 
        \COREAXI_0_AXImslave16_ARSIZE[1]\, 
        \COREAXI_0_AXImslave16_ARBURST[0]\, \axi_state[6]\, 
        \RDATA_reg[46]\, \RDATA_reg[43]\, 
        \COREAXI_0_AXImslave16_RDATA[14]\, 
        \COREAXI_0_AXImslave16_RDATA[11]\, 
        \COREAXI_0_AXImslave16_RDATA_m[57]\, 
        \COREAXI_0_AXImslave16_RDATA_m[58]\, 
        \COREAXI_0_AXImslave16_RDATA_m[41]\, 
        \COREAXI_0_AXImslave16_RDATA_m[42]\, 
        \COREAXI_0_AXImslave16_RDATA_m[47]\, 
        \COREAXI_0_AXImslave16_RDATA_m[49]\, 
        \COREAXI_0_AXImslave16_RDATA_m[50]\, 
        \COREAXI_0_AXImslave16_RDATA_m[33]\, 
        \COREAXI_0_AXImslave16_RDATA_m[34]\, 
        \COREAXI_0_AXImslave16_RDATA_m[11]\, 
        \COREAXI_0_AXImslave16_RDATA_m[12]\, 
        \COREAXI_0_AXImslave16_RDATA_m[13]\, 
        \COREAXI_0_AXImslave16_RDATA_m[14]\, 
        \COREAXI_0_AXImslave16_RDATA_m[15]\, 
        \COREAXI_0_AXImslave16_RDATA_m[19]\, 
        \COREAXI_0_AXImslave16_RDATA_m[20]\, 
        \COREAXI_0_AXImslave16_RDATA_m[21]\, 
        \COREAXI_0_AXImslave16_RDATA_m[23]\, 
        \COREAXI_0_AXImslave16_RDATA_m[0]\, 
        \COREAXI_0_AXImslave16_RDATA_m[1]\, 
        \COREAXI_0_AXImslave16_RDATA_m[4]\, 
        \COREAXI_0_AXImslave16_RDATA_m[5]\, 
        \COREAXI_0_AXImslave16_RDATA_m[6]\, 
        \COREAXI_0_AXImslave16_RDATA_m[7]\, 
        \COREAXI_0_AXImslave16_RDATA_m[8]\, 
        \COREAXI_0_AXImslave16_RDATA_m[9]\, 
        \COREAXI_0_AXImslave16_RDATA_m[10]\, 
        COREAXI_0_AXImslave16_WVALID, WREADY_SI16_i, 
        COREAXI_0_AXImslave16_AWVALID, 
        COREAXI_0_AXImslave16_AWREADY, 
        COREAXI_0_AXImslave16_BVALID, N_3297, N_389, N_74, 
        N_3167_i, N_23, N_3170_i, N_39, N_78_mux_i, N_79_mux_i, 
        N_80_mux_i, N_70_mux_i, N_71_mux_i, N_72_mux_i, N_3094_i, 
        N_3096_i, N_3098_i, N_3100_i, N_3102_i, N_3169_i, 
        N_3066_i, N_67_mux_i, N_68_mux_i, N_69_mux_i, N_75_mux_i, 
        N_76_mux_i, N_77_mux_i, i22_mux_2_i, i22_mux_3_i, 
        i22_mux_4_i, i22_mux_5_i, N_8_i, i17_mux_2_i, N_3064_i, 
        N_3092_i, i17_mux_i, i17_mux_0_i, i17_mux_1_i, i22_mux_i, 
        i22_mux_0_i, i22_mux_1_i, COREAXI_0_AXImslave16_ARREADY, 
        COREAXI_0_AXImslave16_ARVALID, WREADY_SI16, 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        top_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CORERESETP_0_RESET_N_F2M, GND_net_1, VCC_net_1
         : std_logic;
    signal nc10, nc8, nc7, nc6, nc2, nc9, nc5, nc4, nc3, nc1
         : std_logic;

    for all : CORESDR_AXI
	Use entity work.CORESDR_AXI(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : CoreAHBLite
	Use entity work.CoreAHBLite(DEF_ARCH);
    for all : top_sb_CCC_0_FCCC
	Use entity work.top_sb_CCC_0_FCCC(DEF_ARCH);
    for all : top_sb_MSS
	Use entity work.top_sb_MSS(DEF_ARCH);
    for all : top_sb_COREAXI_0_COREAXI
	Use entity work.top_sb_COREAXI_0_COREAXI(DEF_ARCH);
    for all : top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI
	Use entity work.top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI(DEF_ARCH);
begin 

    SDRCLK_c <= \SDRCLK_c\;

    MSS_SMC_0 : CORESDR_AXI
      port map(COREAXI_0_AXImslave16_AWSIZE(1) => 
        \COREAXI_0_AXImslave16_AWSIZE[1]\, 
        COREAXI_0_AXImslave16_AWSIZE(0) => 
        \COREAXI_0_AXImslave16_AWSIZE[0]\, 
        COREAXI_0_AXImslave16_ARSIZE(1) => 
        \COREAXI_0_AXImslave16_ARSIZE[1]\, 
        COREAXI_0_AXImslave16_ARSIZE(0) => 
        \COREAXI_0_AXImslave16_ARSIZE[0]\, 
        COREAXI_0_AXImslave16_WDATA(63) => 
        \COREAXI_0_AXImslave16_WDATA[63]\, 
        COREAXI_0_AXImslave16_WDATA(62) => 
        \COREAXI_0_AXImslave16_WDATA[62]\, 
        COREAXI_0_AXImslave16_WDATA(61) => 
        \COREAXI_0_AXImslave16_WDATA[61]\, 
        COREAXI_0_AXImslave16_WDATA(60) => 
        \COREAXI_0_AXImslave16_WDATA[60]\, 
        COREAXI_0_AXImslave16_WDATA(59) => 
        \COREAXI_0_AXImslave16_WDATA[59]\, 
        COREAXI_0_AXImslave16_WDATA(58) => 
        \COREAXI_0_AXImslave16_WDATA[58]\, 
        COREAXI_0_AXImslave16_WDATA(57) => 
        \COREAXI_0_AXImslave16_WDATA[57]\, 
        COREAXI_0_AXImslave16_WDATA(56) => 
        \COREAXI_0_AXImslave16_WDATA[56]\, 
        COREAXI_0_AXImslave16_WDATA(55) => 
        \COREAXI_0_AXImslave16_WDATA[55]\, 
        COREAXI_0_AXImslave16_WDATA(54) => 
        \COREAXI_0_AXImslave16_WDATA[54]\, 
        COREAXI_0_AXImslave16_WDATA(53) => 
        \COREAXI_0_AXImslave16_WDATA[53]\, 
        COREAXI_0_AXImslave16_WDATA(52) => 
        \COREAXI_0_AXImslave16_WDATA[52]\, 
        COREAXI_0_AXImslave16_WDATA(51) => 
        \COREAXI_0_AXImslave16_WDATA[51]\, 
        COREAXI_0_AXImslave16_WDATA(50) => 
        \COREAXI_0_AXImslave16_WDATA[50]\, 
        COREAXI_0_AXImslave16_WDATA(49) => 
        \COREAXI_0_AXImslave16_WDATA[49]\, 
        COREAXI_0_AXImslave16_WDATA(48) => 
        \COREAXI_0_AXImslave16_WDATA[48]\, 
        COREAXI_0_AXImslave16_WDATA(47) => 
        \COREAXI_0_AXImslave16_WDATA[47]\, 
        COREAXI_0_AXImslave16_WDATA(46) => 
        \COREAXI_0_AXImslave16_WDATA[46]\, 
        COREAXI_0_AXImslave16_WDATA(45) => 
        \COREAXI_0_AXImslave16_WDATA[45]\, 
        COREAXI_0_AXImslave16_WDATA(44) => 
        \COREAXI_0_AXImslave16_WDATA[44]\, 
        COREAXI_0_AXImslave16_WDATA(43) => 
        \COREAXI_0_AXImslave16_WDATA[43]\, 
        COREAXI_0_AXImslave16_WDATA(42) => 
        \COREAXI_0_AXImslave16_WDATA[42]\, 
        COREAXI_0_AXImslave16_WDATA(41) => 
        \COREAXI_0_AXImslave16_WDATA[41]\, 
        COREAXI_0_AXImslave16_WDATA(40) => 
        \COREAXI_0_AXImslave16_WDATA[40]\, 
        COREAXI_0_AXImslave16_WDATA(39) => 
        \COREAXI_0_AXImslave16_WDATA[39]\, 
        COREAXI_0_AXImslave16_WDATA(38) => 
        \COREAXI_0_AXImslave16_WDATA[38]\, 
        COREAXI_0_AXImslave16_WDATA(37) => 
        \COREAXI_0_AXImslave16_WDATA[37]\, 
        COREAXI_0_AXImslave16_WDATA(36) => 
        \COREAXI_0_AXImslave16_WDATA[36]\, 
        COREAXI_0_AXImslave16_WDATA(35) => 
        \COREAXI_0_AXImslave16_WDATA[35]\, 
        COREAXI_0_AXImslave16_WDATA(34) => 
        \COREAXI_0_AXImslave16_WDATA[34]\, 
        COREAXI_0_AXImslave16_WDATA(33) => 
        \COREAXI_0_AXImslave16_WDATA[33]\, 
        COREAXI_0_AXImslave16_WDATA(32) => 
        \COREAXI_0_AXImslave16_WDATA[32]\, 
        COREAXI_0_AXImslave16_WDATA(31) => 
        \COREAXI_0_AXImslave16_WDATA[31]\, 
        COREAXI_0_AXImslave16_WDATA(30) => 
        \COREAXI_0_AXImslave16_WDATA[30]\, 
        COREAXI_0_AXImslave16_WDATA(29) => 
        \COREAXI_0_AXImslave16_WDATA[29]\, 
        COREAXI_0_AXImslave16_WDATA(28) => 
        \COREAXI_0_AXImslave16_WDATA[28]\, 
        COREAXI_0_AXImslave16_WDATA(27) => 
        \COREAXI_0_AXImslave16_WDATA[27]\, 
        COREAXI_0_AXImslave16_WDATA(26) => 
        \COREAXI_0_AXImslave16_WDATA[26]\, 
        COREAXI_0_AXImslave16_WDATA(25) => 
        \COREAXI_0_AXImslave16_WDATA[25]\, 
        COREAXI_0_AXImslave16_WDATA(24) => 
        \COREAXI_0_AXImslave16_WDATA[24]\, 
        COREAXI_0_AXImslave16_WDATA(23) => 
        \COREAXI_0_AXImslave16_WDATA[23]\, 
        COREAXI_0_AXImslave16_WDATA(22) => 
        \COREAXI_0_AXImslave16_WDATA[22]\, 
        COREAXI_0_AXImslave16_WDATA(21) => 
        \COREAXI_0_AXImslave16_WDATA[21]\, 
        COREAXI_0_AXImslave16_WDATA(20) => 
        \COREAXI_0_AXImslave16_WDATA[20]\, 
        COREAXI_0_AXImslave16_WDATA(19) => 
        \COREAXI_0_AXImslave16_WDATA[19]\, 
        COREAXI_0_AXImslave16_WDATA(18) => 
        \COREAXI_0_AXImslave16_WDATA[18]\, 
        COREAXI_0_AXImslave16_WDATA(17) => 
        \COREAXI_0_AXImslave16_WDATA[17]\, 
        COREAXI_0_AXImslave16_WDATA(16) => 
        \COREAXI_0_AXImslave16_WDATA[16]\, 
        COREAXI_0_AXImslave16_WDATA(15) => 
        \COREAXI_0_AXImslave16_WDATA[15]\, 
        COREAXI_0_AXImslave16_WDATA(14) => 
        \COREAXI_0_AXImslave16_WDATA[14]\, 
        COREAXI_0_AXImslave16_WDATA(13) => 
        \COREAXI_0_AXImslave16_WDATA[13]\, 
        COREAXI_0_AXImslave16_WDATA(12) => 
        \COREAXI_0_AXImslave16_WDATA[12]\, 
        COREAXI_0_AXImslave16_WDATA(11) => 
        \COREAXI_0_AXImslave16_WDATA[11]\, 
        COREAXI_0_AXImslave16_WDATA(10) => 
        \COREAXI_0_AXImslave16_WDATA[10]\, 
        COREAXI_0_AXImslave16_WDATA(9) => 
        \COREAXI_0_AXImslave16_WDATA[9]\, 
        COREAXI_0_AXImslave16_WDATA(8) => 
        \COREAXI_0_AXImslave16_WDATA[8]\, 
        COREAXI_0_AXImslave16_WDATA(7) => 
        \COREAXI_0_AXImslave16_WDATA[7]\, 
        COREAXI_0_AXImslave16_WDATA(6) => 
        \COREAXI_0_AXImslave16_WDATA[6]\, 
        COREAXI_0_AXImslave16_WDATA(5) => 
        \COREAXI_0_AXImslave16_WDATA[5]\, 
        COREAXI_0_AXImslave16_WDATA(4) => 
        \COREAXI_0_AXImslave16_WDATA[4]\, 
        COREAXI_0_AXImslave16_WDATA(3) => 
        \COREAXI_0_AXImslave16_WDATA[3]\, 
        COREAXI_0_AXImslave16_WDATA(2) => 
        \COREAXI_0_AXImslave16_WDATA[2]\, 
        COREAXI_0_AXImslave16_WDATA(1) => 
        \COREAXI_0_AXImslave16_WDATA[1]\, 
        COREAXI_0_AXImslave16_WDATA(0) => 
        \COREAXI_0_AXImslave16_WDATA[0]\, 
        COREAXI_0_AXImslave16_AWADDR(23) => 
        \COREAXI_0_AXImslave16_AWADDR[23]\, 
        COREAXI_0_AXImslave16_AWADDR(22) => 
        \COREAXI_0_AXImslave16_AWADDR[22]\, 
        COREAXI_0_AXImslave16_AWADDR(21) => 
        \COREAXI_0_AXImslave16_AWADDR[21]\, 
        COREAXI_0_AXImslave16_AWADDR(20) => 
        \COREAXI_0_AXImslave16_AWADDR[20]\, 
        COREAXI_0_AXImslave16_AWADDR(19) => 
        \COREAXI_0_AXImslave16_AWADDR[19]\, 
        COREAXI_0_AXImslave16_AWADDR(18) => 
        \COREAXI_0_AXImslave16_AWADDR[18]\, 
        COREAXI_0_AXImslave16_AWADDR(17) => 
        \COREAXI_0_AXImslave16_AWADDR[17]\, 
        COREAXI_0_AXImslave16_AWADDR(16) => 
        \COREAXI_0_AXImslave16_AWADDR[16]\, 
        COREAXI_0_AXImslave16_AWADDR(15) => 
        \COREAXI_0_AXImslave16_AWADDR[15]\, 
        COREAXI_0_AXImslave16_AWADDR(14) => 
        \COREAXI_0_AXImslave16_AWADDR[14]\, 
        COREAXI_0_AXImslave16_AWADDR(13) => 
        \COREAXI_0_AXImslave16_AWADDR[13]\, 
        COREAXI_0_AXImslave16_AWADDR(12) => 
        \COREAXI_0_AXImslave16_AWADDR[12]\, 
        COREAXI_0_AXImslave16_AWADDR(11) => 
        \COREAXI_0_AXImslave16_AWADDR[11]\, 
        COREAXI_0_AXImslave16_AWADDR(10) => 
        \COREAXI_0_AXImslave16_AWADDR[10]\, 
        COREAXI_0_AXImslave16_AWADDR(9) => 
        \COREAXI_0_AXImslave16_AWADDR[9]\, 
        COREAXI_0_AXImslave16_AWADDR(8) => 
        \COREAXI_0_AXImslave16_AWADDR[8]\, 
        COREAXI_0_AXImslave16_AWADDR(7) => 
        \COREAXI_0_AXImslave16_AWADDR[7]\, 
        COREAXI_0_AXImslave16_AWADDR(6) => 
        \COREAXI_0_AXImslave16_AWADDR[6]\, 
        COREAXI_0_AXImslave16_AWADDR(5) => 
        \COREAXI_0_AXImslave16_AWADDR[5]\, 
        COREAXI_0_AXImslave16_AWADDR(4) => 
        \COREAXI_0_AXImslave16_AWADDR[4]\, 
        COREAXI_0_AXImslave16_AWADDR(3) => 
        \COREAXI_0_AXImslave16_AWADDR[3]\, 
        COREAXI_0_AXImslave16_AWADDR(2) => 
        \COREAXI_0_AXImslave16_AWADDR[2]\, 
        COREAXI_0_AXImslave16_AWADDR(1) => 
        \COREAXI_0_AXImslave16_AWADDR[1]\, 
        COREAXI_0_AXImslave16_ARADDR(23) => 
        \COREAXI_0_AXImslave16_ARADDR[23]\, 
        COREAXI_0_AXImslave16_ARADDR(22) => 
        \COREAXI_0_AXImslave16_ARADDR[22]\, 
        COREAXI_0_AXImslave16_ARADDR(21) => 
        \COREAXI_0_AXImslave16_ARADDR[21]\, 
        COREAXI_0_AXImslave16_ARADDR(20) => 
        \COREAXI_0_AXImslave16_ARADDR[20]\, 
        COREAXI_0_AXImslave16_ARADDR(19) => 
        \COREAXI_0_AXImslave16_ARADDR[19]\, 
        COREAXI_0_AXImslave16_ARADDR(18) => 
        \COREAXI_0_AXImslave16_ARADDR[18]\, 
        COREAXI_0_AXImslave16_ARADDR(17) => 
        \COREAXI_0_AXImslave16_ARADDR[17]\, 
        COREAXI_0_AXImslave16_ARADDR(16) => 
        \COREAXI_0_AXImslave16_ARADDR[16]\, 
        COREAXI_0_AXImslave16_ARADDR(15) => 
        \COREAXI_0_AXImslave16_ARADDR[15]\, 
        COREAXI_0_AXImslave16_ARADDR(14) => 
        \COREAXI_0_AXImslave16_ARADDR[14]\, 
        COREAXI_0_AXImslave16_ARADDR(13) => 
        \COREAXI_0_AXImslave16_ARADDR[13]\, 
        COREAXI_0_AXImslave16_ARADDR(12) => 
        \COREAXI_0_AXImslave16_ARADDR[12]\, 
        COREAXI_0_AXImslave16_ARADDR(11) => 
        \COREAXI_0_AXImslave16_ARADDR[11]\, 
        COREAXI_0_AXImslave16_ARADDR(10) => 
        \COREAXI_0_AXImslave16_ARADDR[10]\, 
        COREAXI_0_AXImslave16_ARADDR(9) => 
        \COREAXI_0_AXImslave16_ARADDR[9]\, 
        COREAXI_0_AXImslave16_ARADDR(8) => 
        \COREAXI_0_AXImslave16_ARADDR[8]\, 
        COREAXI_0_AXImslave16_ARADDR(7) => 
        \COREAXI_0_AXImslave16_ARADDR[7]\, 
        COREAXI_0_AXImslave16_ARADDR(6) => 
        \COREAXI_0_AXImslave16_ARADDR[6]\, 
        COREAXI_0_AXImslave16_ARADDR(5) => 
        \COREAXI_0_AXImslave16_ARADDR[5]\, 
        COREAXI_0_AXImslave16_ARADDR(4) => 
        \COREAXI_0_AXImslave16_ARADDR[4]\, 
        COREAXI_0_AXImslave16_ARADDR(3) => 
        \COREAXI_0_AXImslave16_ARADDR[3]\, 
        COREAXI_0_AXImslave16_ARADDR(2) => 
        \COREAXI_0_AXImslave16_ARADDR[2]\, 
        COREAXI_0_AXImslave16_ARADDR(1) => 
        \COREAXI_0_AXImslave16_ARADDR[1]\, 
        COREAXI_0_AXImslave16_WSTRB(7) => 
        \COREAXI_0_AXImslave16_WSTRB[7]\, 
        COREAXI_0_AXImslave16_WSTRB(6) => 
        \COREAXI_0_AXImslave16_WSTRB[6]\, 
        COREAXI_0_AXImslave16_WSTRB(5) => 
        \COREAXI_0_AXImslave16_WSTRB[5]\, 
        COREAXI_0_AXImslave16_WSTRB(4) => 
        \COREAXI_0_AXImslave16_WSTRB[4]\, 
        COREAXI_0_AXImslave16_WSTRB(3) => 
        \COREAXI_0_AXImslave16_WSTRB[3]\, 
        COREAXI_0_AXImslave16_WSTRB(2) => 
        \COREAXI_0_AXImslave16_WSTRB[2]\, 
        COREAXI_0_AXImslave16_WSTRB(1) => 
        \COREAXI_0_AXImslave16_WSTRB[1]\, 
        COREAXI_0_AXImslave16_WSTRB(0) => 
        \COREAXI_0_AXImslave16_WSTRB[0]\, DQM_c(1) => DQM_c(1), 
        DQM_c(0) => DQM_c(0), sdr_datain_reg(15) => 
        sdr_datain_reg(15), sdr_datain_reg(14) => 
        sdr_datain_reg(14), sdr_datain_reg(13) => 
        sdr_datain_reg(13), sdr_datain_reg(12) => 
        sdr_datain_reg(12), sdr_datain_reg(11) => 
        sdr_datain_reg(11), sdr_datain_reg(10) => 
        sdr_datain_reg(10), sdr_datain_reg(9) => 
        sdr_datain_reg(9), sdr_datain_reg(8) => sdr_datain_reg(8), 
        sdr_datain_reg(7) => sdr_datain_reg(7), sdr_datain_reg(6)
         => sdr_datain_reg(6), sdr_datain_reg(5) => 
        sdr_datain_reg(5), sdr_datain_reg(4) => sdr_datain_reg(4), 
        sdr_datain_reg(3) => sdr_datain_reg(3), sdr_datain_reg(2)
         => sdr_datain_reg(2), sdr_datain_reg(1) => 
        sdr_datain_reg(1), sdr_datain_reg(0) => sdr_datain_reg(0), 
        SA_c(11) => SA_c(11), SA_c(10) => SA_c(10), SA_c(9) => 
        SA_c(9), SA_c(8) => SA_c(8), SA_c(7) => SA_c(7), SA_c(6)
         => SA_c(6), SA_c(5) => SA_c(5), SA_c(4) => SA_c(4), 
        SA_c(3) => SA_c(3), SA_c(2) => SA_c(2), SA_c(1) => 
        SA_c(1), SA_c(0) => SA_c(0), BA_c(1) => BA_c(1), BA_c(0)
         => BA_c(0), DQ_in(15) => DQ_in(15), DQ_in(14) => 
        DQ_in(14), DQ_in(13) => DQ_in(13), DQ_in(12) => DQ_in(12), 
        DQ_in(11) => DQ_in(11), DQ_in(10) => DQ_in(10), DQ_in(9)
         => DQ_in(9), DQ_in(8) => DQ_in(8), DQ_in(7) => DQ_in(7), 
        DQ_in(6) => DQ_in(6), DQ_in(5) => DQ_in(5), DQ_in(4) => 
        DQ_in(4), DQ_in(3) => DQ_in(3), DQ_in(2) => DQ_in(2), 
        DQ_in(1) => DQ_in(1), DQ_in(0) => DQ_in(0), 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        \COREAXI_0_AXImslave16_RDATA_m[8]\, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        \COREAXI_0_AXImslave16_RDATA_m[11]\, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        \COREAXI_0_AXImslave16_RDATA_m[12]\, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        \COREAXI_0_AXImslave16_RDATA_m[13]\, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        \COREAXI_0_AXImslave16_RDATA_m[14]\, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        \COREAXI_0_AXImslave16_RDATA_m[15]\, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        \COREAXI_0_AXImslave16_RDATA_m[0]\, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        \COREAXI_0_AXImslave16_RDATA_m[4]\, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        \COREAXI_0_AXImslave16_RDATA_m[5]\, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        \COREAXI_0_AXImslave16_RDATA_m[6]\, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        \COREAXI_0_AXImslave16_RDATA_m[7]\, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        \COREAXI_0_AXImslave16_RDATA_m[10]\, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        \COREAXI_0_AXImslave16_RDATA_m[9]\, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        \COREAXI_0_AXImslave16_RDATA_m[1]\, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        \COREAXI_0_AXImslave16_RDATA_m[34]\, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        \COREAXI_0_AXImslave16_RDATA_m[47]\, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        \COREAXI_0_AXImslave16_RDATA_m[19]\, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        \COREAXI_0_AXImslave16_RDATA_m[20]\, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        \COREAXI_0_AXImslave16_RDATA_m[21]\, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        \COREAXI_0_AXImslave16_RDATA_m[23]\, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        \COREAXI_0_AXImslave16_RDATA_m[41]\, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        \COREAXI_0_AXImslave16_RDATA_m[33]\, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        \COREAXI_0_AXImslave16_RDATA_m[42]\, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        \COREAXI_0_AXImslave16_RDATA_m[49]\, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        \COREAXI_0_AXImslave16_RDATA_m[50]\, 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        \COREAXI_0_AXImslave16_RDATA_m[57]\, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        \COREAXI_0_AXImslave16_RDATA_m[58]\, 
        COREAXI_0_AXImslave16_ARBURST_0 => 
        \COREAXI_0_AXImslave16_ARBURST[0]\, CS_N_c_0 => CS_N_c_0, 
        axi_state_0 => \axi_state[6]\, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        \COREAXI_0_AXImslave16_RDATA[11]\, 
        COREAXI_0_AXImslave16_RDATA_3 => 
        \COREAXI_0_AXImslave16_RDATA[14]\, RDATA_reg_0 => 
        \RDATA_reg[43]\, RDATA_reg_3 => \RDATA_reg[46]\, N_8_i
         => N_8_i, N_23 => N_23, N_3169_i => N_3169_i, N_77_mux_i
         => N_77_mux_i, N_76_mux_i => N_76_mux_i, N_75_mux_i => 
        N_75_mux_i, N_69_mux_i => N_69_mux_i, N_68_mux_i => 
        N_68_mux_i, N_67_mux_i => N_67_mux_i, N_72_mux_i => 
        N_72_mux_i, N_71_mux_i => N_71_mux_i, N_70_mux_i => 
        N_70_mux_i, N_80_mux_i => N_80_mux_i, N_79_mux_i => 
        N_79_mux_i, N_78_mux_i => N_78_mux_i, N_3297 => N_3297, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID, N_3170_i => N_3170_i, 
        COREAXI_0_AXImslave16_AWVALID => 
        COREAXI_0_AXImslave16_AWVALID, N_39 => N_39, 
        WREADY_SI16_i => WREADY_SI16_i, 
        COREAXI_0_AXImslave16_WVALID => 
        COREAXI_0_AXImslave16_WVALID, 
        COREAXI_0_AXImslave16_ARVALID => 
        COREAXI_0_AXImslave16_ARVALID, i22_mux_2_i => i22_mux_2_i, 
        i22_mux_3_i => i22_mux_3_i, i22_mux_4_i => i22_mux_4_i, 
        i22_mux_5_i => i22_mux_5_i, i17_mux_2_i => i17_mux_2_i, 
        i17_mux_i => i17_mux_i, i17_mux_0_i => i17_mux_0_i, 
        i17_mux_1_i => i17_mux_1_i, i22_mux_i => i22_mux_i, 
        i22_mux_0_i => i22_mux_0_i, i22_mux_1_i => i22_mux_1_i, 
        N_389 => N_389, N_3064_i => N_3064_i, N_3066_i => 
        N_3066_i, N_3092_i => N_3092_i, N_3094_i => N_3094_i, 
        N_3096_i => N_3096_i, N_3098_i => N_3098_i, N_3100_i => 
        N_3100_i, N_3102_i => N_3102_i, N_74 => N_74, N_3167_i
         => N_3167_i, WE_N_c => WE_N_c, RAS_N_c => RAS_N_c, 
        un1_top_sb_0_3_i_i => un1_top_sb_0_3_i_i, CKE_c => CKE_c, 
        CAS_N_c => CAS_N_c, COREAXI_0_AXImslave16_BVALID => 
        COREAXI_0_AXImslave16_BVALID, 
        COREAXI_0_AXImslave16_AWREADY => 
        COREAXI_0_AXImslave16_AWREADY, 
        COREAXI_0_AXImslave16_ARREADY => 
        COREAXI_0_AXImslave16_ARREADY, WREADY_SI16 => WREADY_SI16, 
        SDRCLK_c => \SDRCLK_c\, MSS_READY => MSS_READY);
    
    CORERESETP_0 : CoreResetP
      port map(top_sb_0_POWER_ON_RESET_N => 
        top_sb_0_POWER_ON_RESET_N, 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        top_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        top_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CORERESETP_0_RESET_N_F2M => CORERESETP_0_RESET_N_F2M, 
        SDRCLK_c => \SDRCLK_c\, MSS_READY => MSS_READY);
    
    CoreAHBLite_0 : CoreAHBLite
      port map(top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[31]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[30]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[29]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[28]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[27]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[26]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[25]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[24]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[23]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[22]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[21]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[20]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[19]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[18]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[17]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[16]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[15]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[14]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[13]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[12]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[11]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[9]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[8]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[7]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[6]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[5]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[4]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[3]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[2]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[0]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(27) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[27]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(26) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[26]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(25) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[25]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(24) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[24]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(23) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[23]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(22) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[22]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(21) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[21]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(20) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[20]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(19) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[19]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(18) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[18]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(17) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[17]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(16) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[16]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(15) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[15]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(14) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[14]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(13) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[13]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(12) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[12]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(11) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[11]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(10) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[10]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(9) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[9]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(8) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[8]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(7) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[7]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(6) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[6]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(5) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[5]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(4) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[4]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(3) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[3]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(2) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[2]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(1) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[1]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(0) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[0]\, 
        CoreAHBLite_0_AHBmslave10_HSIZE(1) => 
        \CoreAHBLite_0_AHBmslave10_HSIZE[1]\, 
        CoreAHBLite_0_AHBmslave10_HSIZE(0) => 
        \CoreAHBLite_0_AHBmslave10_HSIZE[0]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(31) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[31]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(30) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[30]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(29) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[29]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(28) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[28]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(27) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[27]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(26) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[26]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(25) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[25]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(24) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[24]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(23) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[23]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(22) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[22]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(21) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[21]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(20) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[20]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(19) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[19]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(18) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[18]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(17) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[17]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(16) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[16]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(15) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[15]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(14) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[14]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(13) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[13]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(12) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[12]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(11) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[11]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(10) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[10]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(9) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[9]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(8) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[8]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(7) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[7]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(6) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[6]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(5) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[5]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(4) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[4]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(3) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[3]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(2) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[2]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(1) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[1]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(0) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[31]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[30]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[29]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[28]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[27]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[26]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[25]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[24]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[23]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[22]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[21]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[20]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[19]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[18]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[17]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[16]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[15]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[14]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[13]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[12]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[11]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[9]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[8]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[7]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[6]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[5]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[4]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[3]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[2]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[0]\, 
        masterAddrInProg_0 => \masterAddrInProg[0]\, 
        current_state_0 => \current_state[7]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0 => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP[0]\, 
        xhdl1222_0 => \xhdl1222[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY, N_92 => N_92, 
        N_91 => N_91, hready_m_xhdl349 => hready_m_xhdl349, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        m0PrevDataSlaveReady => m0PrevDataSlaveReady, SDRCLK_c
         => \SDRCLK_c\, MSS_READY => MSS_READY, 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK => 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, 
        CoreAHBLite_0_AHBmslave10_HWRITE => 
        CoreAHBLite_0_AHBmslave10_HWRITE, hsel2 => hsel2, 
        hsel2_0_a2_1 => hsel2_0_a2_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CCC_0 : top_sb_CCC_0_FCCC
      port map(FAB_CCC_LOCK => FAB_CCC_LOCK, CLK1_PAD => CLK1_PAD, 
        SDRCLK_c => \SDRCLK_c\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    top_sb_MSS_0 : top_sb_MSS
      port map(top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HSIZE[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(31) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[31]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(30) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[30]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(29) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[29]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(28) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[28]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(27) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[27]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(26) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[26]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(25) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[25]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(24) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[24]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(23) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[23]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(22) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[22]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(21) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[21]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(20) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[20]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(19) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[19]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(18) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[18]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(17) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[17]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(16) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[16]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(15) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[15]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(14) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[14]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(13) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[13]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(12) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[12]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(11) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[11]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(10) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(9) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[9]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(8) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[8]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(7) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[7]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(6) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[6]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(5) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[5]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(4) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[4]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(3) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[3]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(2) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[2]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWDATA[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(31) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[31]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(30) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[30]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(29) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[29]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(28) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[28]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(27) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[27]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(26) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[26]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(25) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[25]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(24) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[24]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(23) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[23]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(22) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[22]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(21) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[21]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(20) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[20]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(19) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[19]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(18) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[18]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(17) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[17]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(16) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[16]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(15) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[15]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(14) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[14]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(13) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[13]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(12) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[12]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(11) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[11]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(10) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[10]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(9) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[9]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(8) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[8]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(7) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[7]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(6) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[6]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(5) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[5]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(4) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[4]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(3) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[3]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(2) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[2]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(1) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR(0) => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HADDR[0]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP_0 => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HRESP[0]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS_0 => 
        \top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HTRANS[1]\, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HREADY, SDRCLK_c => 
        \SDRCLK_c\, CORERESETP_0_RESET_N_F2M => 
        CORERESETP_0_RESET_N_F2M, FAB_CCC_LOCK => FAB_CCC_LOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HLOCK, 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE => 
        top_sb_MSS_TMP_0_MDDR_SMC_AHB_MASTER_HWRITE, 
        top_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        top_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N => 
        top_sb_MSS_TMP_0_FIC_2_APB_M_PRESET_N, hready_m_xhdl349
         => hready_m_xhdl349, CAN_RX => CAN_RX, CAN_TX_EN_N => 
        CAN_TX_EN_N, CAN_TX => CAN_TX, GPIO_1_BI => GPIO_1_BI, 
        GPIO_8_BI => GPIO_8_BI, GPIO_9_BI => GPIO_9_BI, 
        GPIO_10_BI => GPIO_10_BI, GPIO_11_BI => GPIO_11_BI, 
        GPIO_12_BI => GPIO_12_BI, GPIO_13_BI => GPIO_13_BI, 
        GPIO_14_BI => GPIO_14_BI, GPIO_15_BI => GPIO_15_BI, 
        GPIO_16_BI => GPIO_16_BI, GPIO_17_BI => GPIO_17_BI, 
        GPIO_18_BI => GPIO_18_BI, GPIO_19_BI => GPIO_19_BI, 
        GPIO_20_BI => GPIO_20_BI, GPIO_21_BI => GPIO_21_BI, 
        GPIO_22_BI => GPIO_22_BI, GPIO_23_BI => GPIO_23_BI, 
        GPIO_24_BI => GPIO_24_BI, GPIO_25_BI => GPIO_25_BI, 
        GPIO_26_BI => GPIO_26_BI, GPIO_29_BI => GPIO_29_BI, 
        I2C_0_SCL => I2C_0_SCL, I2C_0_SDA => I2C_0_SDA, 
        MMUART_0_RXD => MMUART_0_RXD, MMUART_0_TXD => 
        MMUART_0_TXD, SPI_0_CLK => SPI_0_CLK, SPI_0_DI => 
        SPI_0_DI, SPI_0_DO => SPI_0_DO, SPI_0_SS0 => SPI_0_SS0);
    
    COREAXI_0 : top_sb_COREAXI_0_COREAXI
      port map(COREAXI_0_AXImslave16_AWSIZE(1) => 
        \COREAXI_0_AXImslave16_AWSIZE[1]\, 
        COREAXI_0_AXImslave16_AWSIZE(0) => 
        \COREAXI_0_AXImslave16_AWSIZE[0]\, 
        COREAXI_0_AXImslave16_ARADDR(23) => 
        \COREAXI_0_AXImslave16_ARADDR[23]\, 
        COREAXI_0_AXImslave16_ARADDR(22) => 
        \COREAXI_0_AXImslave16_ARADDR[22]\, 
        COREAXI_0_AXImslave16_ARADDR(21) => 
        \COREAXI_0_AXImslave16_ARADDR[21]\, 
        COREAXI_0_AXImslave16_ARADDR(20) => 
        \COREAXI_0_AXImslave16_ARADDR[20]\, 
        COREAXI_0_AXImslave16_ARADDR(19) => 
        \COREAXI_0_AXImslave16_ARADDR[19]\, 
        COREAXI_0_AXImslave16_ARADDR(18) => 
        \COREAXI_0_AXImslave16_ARADDR[18]\, 
        COREAXI_0_AXImslave16_ARADDR(17) => 
        \COREAXI_0_AXImslave16_ARADDR[17]\, 
        COREAXI_0_AXImslave16_ARADDR(16) => 
        \COREAXI_0_AXImslave16_ARADDR[16]\, 
        COREAXI_0_AXImslave16_ARADDR(15) => 
        \COREAXI_0_AXImslave16_ARADDR[15]\, 
        COREAXI_0_AXImslave16_ARADDR(14) => 
        \COREAXI_0_AXImslave16_ARADDR[14]\, 
        COREAXI_0_AXImslave16_ARADDR(13) => 
        \COREAXI_0_AXImslave16_ARADDR[13]\, 
        COREAXI_0_AXImslave16_ARADDR(12) => 
        \COREAXI_0_AXImslave16_ARADDR[12]\, 
        COREAXI_0_AXImslave16_ARADDR(11) => 
        \COREAXI_0_AXImslave16_ARADDR[11]\, 
        COREAXI_0_AXImslave16_ARADDR(10) => 
        \COREAXI_0_AXImslave16_ARADDR[10]\, 
        COREAXI_0_AXImslave16_ARADDR(9) => 
        \COREAXI_0_AXImslave16_ARADDR[9]\, 
        COREAXI_0_AXImslave16_ARADDR(8) => 
        \COREAXI_0_AXImslave16_ARADDR[8]\, 
        COREAXI_0_AXImslave16_ARADDR(7) => 
        \COREAXI_0_AXImslave16_ARADDR[7]\, 
        COREAXI_0_AXImslave16_ARADDR(6) => 
        \COREAXI_0_AXImslave16_ARADDR[6]\, 
        COREAXI_0_AXImslave16_ARADDR(5) => 
        \COREAXI_0_AXImslave16_ARADDR[5]\, 
        COREAXI_0_AXImslave16_ARADDR(4) => 
        \COREAXI_0_AXImslave16_ARADDR[4]\, 
        COREAXI_0_AXImslave16_ARADDR(3) => 
        \COREAXI_0_AXImslave16_ARADDR[3]\, 
        COREAXI_0_AXImslave16_ARADDR(2) => 
        \COREAXI_0_AXImslave16_ARADDR[2]\, 
        COREAXI_0_AXImslave16_ARADDR(1) => 
        \COREAXI_0_AXImslave16_ARADDR[1]\, 
        COREAXI_0_AXImslave16_AWADDR(23) => 
        \COREAXI_0_AXImslave16_AWADDR[23]\, 
        COREAXI_0_AXImslave16_AWADDR(22) => 
        \COREAXI_0_AXImslave16_AWADDR[22]\, 
        COREAXI_0_AXImslave16_AWADDR(21) => 
        \COREAXI_0_AXImslave16_AWADDR[21]\, 
        COREAXI_0_AXImslave16_AWADDR(20) => 
        \COREAXI_0_AXImslave16_AWADDR[20]\, 
        COREAXI_0_AXImslave16_AWADDR(19) => 
        \COREAXI_0_AXImslave16_AWADDR[19]\, 
        COREAXI_0_AXImslave16_AWADDR(18) => 
        \COREAXI_0_AXImslave16_AWADDR[18]\, 
        COREAXI_0_AXImslave16_AWADDR(17) => 
        \COREAXI_0_AXImslave16_AWADDR[17]\, 
        COREAXI_0_AXImslave16_AWADDR(16) => 
        \COREAXI_0_AXImslave16_AWADDR[16]\, 
        COREAXI_0_AXImslave16_AWADDR(15) => 
        \COREAXI_0_AXImslave16_AWADDR[15]\, 
        COREAXI_0_AXImslave16_AWADDR(14) => 
        \COREAXI_0_AXImslave16_AWADDR[14]\, 
        COREAXI_0_AXImslave16_AWADDR(13) => 
        \COREAXI_0_AXImslave16_AWADDR[13]\, 
        COREAXI_0_AXImslave16_AWADDR(12) => 
        \COREAXI_0_AXImslave16_AWADDR[12]\, 
        COREAXI_0_AXImslave16_AWADDR(11) => 
        \COREAXI_0_AXImslave16_AWADDR[11]\, 
        COREAXI_0_AXImslave16_AWADDR(10) => 
        \COREAXI_0_AXImslave16_AWADDR[10]\, 
        COREAXI_0_AXImslave16_AWADDR(9) => 
        \COREAXI_0_AXImslave16_AWADDR[9]\, 
        COREAXI_0_AXImslave16_AWADDR(8) => 
        \COREAXI_0_AXImslave16_AWADDR[8]\, 
        COREAXI_0_AXImslave16_AWADDR(7) => 
        \COREAXI_0_AXImslave16_AWADDR[7]\, 
        COREAXI_0_AXImslave16_AWADDR(6) => 
        \COREAXI_0_AXImslave16_AWADDR[6]\, 
        COREAXI_0_AXImslave16_AWADDR(5) => 
        \COREAXI_0_AXImslave16_AWADDR[5]\, 
        COREAXI_0_AXImslave16_AWADDR(4) => 
        \COREAXI_0_AXImslave16_AWADDR[4]\, 
        COREAXI_0_AXImslave16_AWADDR(3) => 
        \COREAXI_0_AXImslave16_AWADDR[3]\, 
        COREAXI_0_AXImslave16_AWADDR(2) => 
        \COREAXI_0_AXImslave16_AWADDR[2]\, 
        COREAXI_0_AXImslave16_AWADDR(1) => 
        \COREAXI_0_AXImslave16_AWADDR[1]\, 
        COREAXI_0_AXImslave16_WSTRB(7) => 
        \COREAXI_0_AXImslave16_WSTRB[7]\, 
        COREAXI_0_AXImslave16_WSTRB(6) => 
        \COREAXI_0_AXImslave16_WSTRB[6]\, 
        COREAXI_0_AXImslave16_WSTRB(5) => 
        \COREAXI_0_AXImslave16_WSTRB[5]\, 
        COREAXI_0_AXImslave16_WSTRB(4) => 
        \COREAXI_0_AXImslave16_WSTRB[4]\, 
        COREAXI_0_AXImslave16_WSTRB(3) => 
        \COREAXI_0_AXImslave16_WSTRB[3]\, 
        COREAXI_0_AXImslave16_WSTRB(2) => 
        \COREAXI_0_AXImslave16_WSTRB[2]\, 
        COREAXI_0_AXImslave16_WSTRB(1) => 
        \COREAXI_0_AXImslave16_WSTRB[1]\, 
        COREAXI_0_AXImslave16_WSTRB(0) => 
        \COREAXI_0_AXImslave16_WSTRB[0]\, 
        COREAXI_0_AXImslave16_WDATA(63) => 
        \COREAXI_0_AXImslave16_WDATA[63]\, 
        COREAXI_0_AXImslave16_WDATA(62) => 
        \COREAXI_0_AXImslave16_WDATA[62]\, 
        COREAXI_0_AXImslave16_WDATA(61) => 
        \COREAXI_0_AXImslave16_WDATA[61]\, 
        COREAXI_0_AXImslave16_WDATA(60) => 
        \COREAXI_0_AXImslave16_WDATA[60]\, 
        COREAXI_0_AXImslave16_WDATA(59) => 
        \COREAXI_0_AXImslave16_WDATA[59]\, 
        COREAXI_0_AXImslave16_WDATA(58) => 
        \COREAXI_0_AXImslave16_WDATA[58]\, 
        COREAXI_0_AXImslave16_WDATA(57) => 
        \COREAXI_0_AXImslave16_WDATA[57]\, 
        COREAXI_0_AXImslave16_WDATA(56) => 
        \COREAXI_0_AXImslave16_WDATA[56]\, 
        COREAXI_0_AXImslave16_WDATA(55) => 
        \COREAXI_0_AXImslave16_WDATA[55]\, 
        COREAXI_0_AXImslave16_WDATA(54) => 
        \COREAXI_0_AXImslave16_WDATA[54]\, 
        COREAXI_0_AXImslave16_WDATA(53) => 
        \COREAXI_0_AXImslave16_WDATA[53]\, 
        COREAXI_0_AXImslave16_WDATA(52) => 
        \COREAXI_0_AXImslave16_WDATA[52]\, 
        COREAXI_0_AXImslave16_WDATA(51) => 
        \COREAXI_0_AXImslave16_WDATA[51]\, 
        COREAXI_0_AXImslave16_WDATA(50) => 
        \COREAXI_0_AXImslave16_WDATA[50]\, 
        COREAXI_0_AXImslave16_WDATA(49) => 
        \COREAXI_0_AXImslave16_WDATA[49]\, 
        COREAXI_0_AXImslave16_WDATA(48) => 
        \COREAXI_0_AXImslave16_WDATA[48]\, 
        COREAXI_0_AXImslave16_WDATA(47) => 
        \COREAXI_0_AXImslave16_WDATA[47]\, 
        COREAXI_0_AXImslave16_WDATA(46) => 
        \COREAXI_0_AXImslave16_WDATA[46]\, 
        COREAXI_0_AXImslave16_WDATA(45) => 
        \COREAXI_0_AXImslave16_WDATA[45]\, 
        COREAXI_0_AXImslave16_WDATA(44) => 
        \COREAXI_0_AXImslave16_WDATA[44]\, 
        COREAXI_0_AXImslave16_WDATA(43) => 
        \COREAXI_0_AXImslave16_WDATA[43]\, 
        COREAXI_0_AXImslave16_WDATA(42) => 
        \COREAXI_0_AXImslave16_WDATA[42]\, 
        COREAXI_0_AXImslave16_WDATA(41) => 
        \COREAXI_0_AXImslave16_WDATA[41]\, 
        COREAXI_0_AXImslave16_WDATA(40) => 
        \COREAXI_0_AXImslave16_WDATA[40]\, 
        COREAXI_0_AXImslave16_WDATA(39) => 
        \COREAXI_0_AXImslave16_WDATA[39]\, 
        COREAXI_0_AXImslave16_WDATA(38) => 
        \COREAXI_0_AXImslave16_WDATA[38]\, 
        COREAXI_0_AXImslave16_WDATA(37) => 
        \COREAXI_0_AXImslave16_WDATA[37]\, 
        COREAXI_0_AXImslave16_WDATA(36) => 
        \COREAXI_0_AXImslave16_WDATA[36]\, 
        COREAXI_0_AXImslave16_WDATA(35) => 
        \COREAXI_0_AXImslave16_WDATA[35]\, 
        COREAXI_0_AXImslave16_WDATA(34) => 
        \COREAXI_0_AXImslave16_WDATA[34]\, 
        COREAXI_0_AXImslave16_WDATA(33) => 
        \COREAXI_0_AXImslave16_WDATA[33]\, 
        COREAXI_0_AXImslave16_WDATA(32) => 
        \COREAXI_0_AXImslave16_WDATA[32]\, 
        COREAXI_0_AXImslave16_WDATA(31) => 
        \COREAXI_0_AXImslave16_WDATA[31]\, 
        COREAXI_0_AXImslave16_WDATA(30) => 
        \COREAXI_0_AXImslave16_WDATA[30]\, 
        COREAXI_0_AXImslave16_WDATA(29) => 
        \COREAXI_0_AXImslave16_WDATA[29]\, 
        COREAXI_0_AXImslave16_WDATA(28) => 
        \COREAXI_0_AXImslave16_WDATA[28]\, 
        COREAXI_0_AXImslave16_WDATA(27) => 
        \COREAXI_0_AXImslave16_WDATA[27]\, 
        COREAXI_0_AXImslave16_WDATA(26) => 
        \COREAXI_0_AXImslave16_WDATA[26]\, 
        COREAXI_0_AXImslave16_WDATA(25) => 
        \COREAXI_0_AXImslave16_WDATA[25]\, 
        COREAXI_0_AXImslave16_WDATA(24) => 
        \COREAXI_0_AXImslave16_WDATA[24]\, 
        COREAXI_0_AXImslave16_WDATA(23) => 
        \COREAXI_0_AXImslave16_WDATA[23]\, 
        COREAXI_0_AXImslave16_WDATA(22) => 
        \COREAXI_0_AXImslave16_WDATA[22]\, 
        COREAXI_0_AXImslave16_WDATA(21) => 
        \COREAXI_0_AXImslave16_WDATA[21]\, 
        COREAXI_0_AXImslave16_WDATA(20) => 
        \COREAXI_0_AXImslave16_WDATA[20]\, 
        COREAXI_0_AXImslave16_WDATA(19) => 
        \COREAXI_0_AXImslave16_WDATA[19]\, 
        COREAXI_0_AXImslave16_WDATA(18) => 
        \COREAXI_0_AXImslave16_WDATA[18]\, 
        COREAXI_0_AXImslave16_WDATA(17) => 
        \COREAXI_0_AXImslave16_WDATA[17]\, 
        COREAXI_0_AXImslave16_WDATA(16) => 
        \COREAXI_0_AXImslave16_WDATA[16]\, 
        COREAXI_0_AXImslave16_WDATA(15) => 
        \COREAXI_0_AXImslave16_WDATA[15]\, 
        COREAXI_0_AXImslave16_WDATA(14) => 
        \COREAXI_0_AXImslave16_WDATA[14]\, 
        COREAXI_0_AXImslave16_WDATA(13) => 
        \COREAXI_0_AXImslave16_WDATA[13]\, 
        COREAXI_0_AXImslave16_WDATA(12) => 
        \COREAXI_0_AXImslave16_WDATA[12]\, 
        COREAXI_0_AXImslave16_WDATA(11) => 
        \COREAXI_0_AXImslave16_WDATA[11]\, 
        COREAXI_0_AXImslave16_WDATA(10) => 
        \COREAXI_0_AXImslave16_WDATA[10]\, 
        COREAXI_0_AXImslave16_WDATA(9) => 
        \COREAXI_0_AXImslave16_WDATA[9]\, 
        COREAXI_0_AXImslave16_WDATA(8) => 
        \COREAXI_0_AXImslave16_WDATA[8]\, 
        COREAXI_0_AXImslave16_WDATA(7) => 
        \COREAXI_0_AXImslave16_WDATA[7]\, 
        COREAXI_0_AXImslave16_WDATA(6) => 
        \COREAXI_0_AXImslave16_WDATA[6]\, 
        COREAXI_0_AXImslave16_WDATA(5) => 
        \COREAXI_0_AXImslave16_WDATA[5]\, 
        COREAXI_0_AXImslave16_WDATA(4) => 
        \COREAXI_0_AXImslave16_WDATA[4]\, 
        COREAXI_0_AXImslave16_WDATA(3) => 
        \COREAXI_0_AXImslave16_WDATA[3]\, 
        COREAXI_0_AXImslave16_WDATA(2) => 
        \COREAXI_0_AXImslave16_WDATA[2]\, 
        COREAXI_0_AXImslave16_WDATA(1) => 
        \COREAXI_0_AXImslave16_WDATA[1]\, 
        COREAXI_0_AXImslave16_WDATA(0) => 
        \COREAXI_0_AXImslave16_WDATA[0]\, 
        COREAXI_0_AXImslave16_ARSIZE(1) => 
        \COREAXI_0_AXImslave16_ARSIZE[1]\, 
        COREAXI_0_AXImslave16_ARSIZE(0) => 
        \COREAXI_0_AXImslave16_ARSIZE[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[63]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[62]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[61]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[60]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[59]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[58]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[57]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[56]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[55]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[54]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[53]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[52]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[51]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[50]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[49]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[48]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[47]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[46]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[45]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[44]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[43]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[42]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[41]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[40]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[39]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[38]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[37]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[36]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[35]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[34]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[33]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[32]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[31]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[30]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[29]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[28]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[21]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[20]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[19]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[16]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[15]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[14]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[13]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[12]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[11]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[10]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[9]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[8]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[7]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[6]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[5]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[4]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[3]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[2]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(63) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[63]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[62]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[61]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[60]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[59]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[58]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[57]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[56]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[55]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[54]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[53]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[52]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[51]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[50]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[49]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[48]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[47]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[46]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[45]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[44]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[43]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[42]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[41]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[40]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[39]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[38]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[37]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[36]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[35]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[34]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[33]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[32]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(31) => nc10, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[30]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[29]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(28) => nc8, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(21) => nc7, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(20) => nc6, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(19) => nc2, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[16]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[21]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[20]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[19]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[16]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[15]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[14]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[13]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[12]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[11]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[10]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[9]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[8]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[7]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[6]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[5]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[4]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[3]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, 
        COREAXI_0_AXImslave16_ARBURST_0 => 
        \COREAXI_0_AXImslave16_ARBURST[0]\, axi_current_state_0
         => \axi_current_state[1]\, axi_current_state_3 => 
        \axi_current_state[4]\, axi_state_0 => \axi_state[6]\, 
        RDATA_reg_3 => \RDATA_reg[46]\, RDATA_reg_0 => 
        \RDATA_reg[43]\, COREAXI_0_AXImslave16_RDATA_3 => 
        \COREAXI_0_AXImslave16_RDATA[14]\, 
        COREAXI_0_AXImslave16_RDATA_0 => 
        \COREAXI_0_AXImslave16_RDATA[11]\, 
        COREAXI_0_AXImslave16_RDATA_m_57 => 
        \COREAXI_0_AXImslave16_RDATA_m[57]\, 
        COREAXI_0_AXImslave16_RDATA_m_58 => 
        \COREAXI_0_AXImslave16_RDATA_m[58]\, 
        COREAXI_0_AXImslave16_RDATA_m_41 => 
        \COREAXI_0_AXImslave16_RDATA_m[41]\, 
        COREAXI_0_AXImslave16_RDATA_m_42 => 
        \COREAXI_0_AXImslave16_RDATA_m[42]\, 
        COREAXI_0_AXImslave16_RDATA_m_47 => 
        \COREAXI_0_AXImslave16_RDATA_m[47]\, 
        COREAXI_0_AXImslave16_RDATA_m_49 => 
        \COREAXI_0_AXImslave16_RDATA_m[49]\, 
        COREAXI_0_AXImslave16_RDATA_m_50 => 
        \COREAXI_0_AXImslave16_RDATA_m[50]\, 
        COREAXI_0_AXImslave16_RDATA_m_33 => 
        \COREAXI_0_AXImslave16_RDATA_m[33]\, 
        COREAXI_0_AXImslave16_RDATA_m_34 => 
        \COREAXI_0_AXImslave16_RDATA_m[34]\, 
        COREAXI_0_AXImslave16_RDATA_m_11 => 
        \COREAXI_0_AXImslave16_RDATA_m[11]\, 
        COREAXI_0_AXImslave16_RDATA_m_12 => 
        \COREAXI_0_AXImslave16_RDATA_m[12]\, 
        COREAXI_0_AXImslave16_RDATA_m_13 => 
        \COREAXI_0_AXImslave16_RDATA_m[13]\, 
        COREAXI_0_AXImslave16_RDATA_m_14 => 
        \COREAXI_0_AXImslave16_RDATA_m[14]\, 
        COREAXI_0_AXImslave16_RDATA_m_15 => 
        \COREAXI_0_AXImslave16_RDATA_m[15]\, 
        COREAXI_0_AXImslave16_RDATA_m_19 => 
        \COREAXI_0_AXImslave16_RDATA_m[19]\, 
        COREAXI_0_AXImslave16_RDATA_m_20 => 
        \COREAXI_0_AXImslave16_RDATA_m[20]\, 
        COREAXI_0_AXImslave16_RDATA_m_21 => 
        \COREAXI_0_AXImslave16_RDATA_m[21]\, 
        COREAXI_0_AXImslave16_RDATA_m_23 => 
        \COREAXI_0_AXImslave16_RDATA_m[23]\, 
        COREAXI_0_AXImslave16_RDATA_m_0 => 
        \COREAXI_0_AXImslave16_RDATA_m[0]\, 
        COREAXI_0_AXImslave16_RDATA_m_1 => 
        \COREAXI_0_AXImslave16_RDATA_m[1]\, 
        COREAXI_0_AXImslave16_RDATA_m_4 => 
        \COREAXI_0_AXImslave16_RDATA_m[4]\, 
        COREAXI_0_AXImslave16_RDATA_m_5 => 
        \COREAXI_0_AXImslave16_RDATA_m[5]\, 
        COREAXI_0_AXImslave16_RDATA_m_6 => 
        \COREAXI_0_AXImslave16_RDATA_m[6]\, 
        COREAXI_0_AXImslave16_RDATA_m_7 => 
        \COREAXI_0_AXImslave16_RDATA_m[7]\, 
        COREAXI_0_AXImslave16_RDATA_m_8 => 
        \COREAXI_0_AXImslave16_RDATA_m[8]\, 
        COREAXI_0_AXImslave16_RDATA_m_9 => 
        \COREAXI_0_AXImslave16_RDATA_m[9]\, 
        COREAXI_0_AXImslave16_RDATA_m_10 => 
        \COREAXI_0_AXImslave16_RDATA_m[10]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARLOCK[1]\, 
        COREAXI_0_AXImslave16_WVALID => 
        COREAXI_0_AXImslave16_WVALID, WREADY_SI16_i => 
        WREADY_SI16_i, COREAXI_0_AXImslave16_AWVALID => 
        COREAXI_0_AXImslave16_AWVALID, 
        COREAXI_0_AXImslave16_AWREADY => 
        COREAXI_0_AXImslave16_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY, wready_m_xhdl2 => 
        wready_m_xhdl2, N_1445_i => N_1445_i, N_1446_i => 
        N_1446_i, N_1447_i => N_1447_i, N_1448_i => N_1448_i, 
        N_1449_i => N_1449_i, N_1450_i => N_1450_i, N_1451_i => 
        N_1451_i, N_1452_i => N_1452_i, N_202_i => N_202_i, 
        N_201_i => N_201_i, N_200_i => N_200_i, N_197_i => 
        N_197_i, N_195_i => N_195_i, N_134_i => N_134_i, N_133_i
         => N_133_i, N_380_i => N_380_i, N_278_i => N_278_i, 
        N_381_i => N_381_i, N_382_i => N_382_i, N_277_i => 
        N_277_i, N_276_i => N_276_i, N_275_i => N_275_i, N_274_i
         => N_274_i, N_273_i => N_273_i, N_272_i => N_272_i, 
        N_203_i => N_203_i, N_137_i => N_137_i, N_136_i => 
        N_136_i, N_135_i => N_135_i, N_48 => N_48, 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_WREADY, araddr_arvalid_clr_d
         => araddr_arvalid_clr_d, 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, awaddr_awvalid_clr_d
         => awaddr_awvalid_clr_d, MSS_READY => MSS_READY, 
        SDRCLK_c => \SDRCLK_c\, COREAXI_0_AXImslave16_BVALID => 
        COREAXI_0_AXImslave16_BVALID, N_3297 => N_3297, N_389 => 
        N_389, N_74 => N_74, N_3167_i => N_3167_i, N_23 => N_23, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, N_3170_i => N_3170_i, 
        N_39 => N_39, N_78_mux_i => N_78_mux_i, N_79_mux_i => 
        N_79_mux_i, N_80_mux_i => N_80_mux_i, N_70_mux_i => 
        N_70_mux_i, N_71_mux_i => N_71_mux_i, N_72_mux_i => 
        N_72_mux_i, N_3094_i => N_3094_i, N_3096_i => N_3096_i, 
        N_3098_i => N_3098_i, N_3100_i => N_3100_i, N_3102_i => 
        N_3102_i, N_3169_i => N_3169_i, N_3066_i => N_3066_i, 
        N_67_mux_i => N_67_mux_i, N_68_mux_i => N_68_mux_i, 
        N_69_mux_i => N_69_mux_i, N_75_mux_i => N_75_mux_i, 
        N_76_mux_i => N_76_mux_i, N_77_mux_i => N_77_mux_i, 
        i22_mux_2_i => i22_mux_2_i, i22_mux_3_i => i22_mux_3_i, 
        i22_mux_4_i => i22_mux_4_i, i22_mux_5_i => i22_mux_5_i, 
        N_8_i => N_8_i, i17_mux_2_i => i17_mux_2_i, N_3064_i => 
        N_3064_i, N_3092_i => N_3092_i, i17_mux_i => i17_mux_i, 
        i17_mux_0_i => i17_mux_0_i, i17_mux_1_i => i17_mux_1_i, 
        i22_mux_i => i22_mux_i, i22_mux_0_i => i22_mux_0_i, 
        i22_mux_1_i => i22_mux_1_i, COREAXI_0_AXImslave16_ARREADY
         => COREAXI_0_AXImslave16_ARREADY, 
        COREAXI_0_AXImslave16_ARVALID => 
        COREAXI_0_AXImslave16_ARVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, WREADY_SI16 => 
        WREADY_SI16, N_75_i => N_75_i);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => top_sb_0_POWER_ON_RESET_N, 
        DEVRST_N => DEVRST_N);
    
    COREAHBLTOAXI_0 : top_sb_COREAHBLTOAXI_0_COREAHBLTOAXI
      port map(COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARSIZE(0) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARSIZE[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(21) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[21]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(20) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[20]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(19) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[19]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[16]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(15) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[15]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(14) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[14]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(13) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[13]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(12) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[12]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(11) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[11]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(10) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[10]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(9) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[9]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(8) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[8]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(7) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[7]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(6) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[6]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(5) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[5]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(4) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[4]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(3) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[3]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(2) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[2]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARADDR(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARADDR[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(63) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[63]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(62) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[62]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(61) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[61]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(60) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[60]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(59) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[59]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(58) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[58]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(57) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[57]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(56) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[56]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(55) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[55]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(54) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[54]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(53) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[53]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(52) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[52]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(51) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[51]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(50) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[50]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(49) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[49]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(48) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[48]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(47) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[47]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(46) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[46]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(45) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[45]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(44) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[44]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(43) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[43]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(42) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[42]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(41) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[41]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(40) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[40]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(39) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[39]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(38) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[38]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(37) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[37]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(36) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[36]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(35) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[35]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(34) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[34]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(33) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[33]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(32) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[32]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(31) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[31]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(30) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[30]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(29) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[29]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(28) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[28]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(21) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[21]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(20) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[20]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(19) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[19]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[16]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(15) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[15]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(14) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[14]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(13) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[13]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(12) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[12]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(11) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[11]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(10) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[10]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(9) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[9]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(8) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[8]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(7) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[7]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(6) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[6]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(5) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[5]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(4) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[4]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(3) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[3]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(2) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[2]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(1) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[1]\, 
        COREAHBLTOAXI_0_AXIMasterIF_RDATA(0) => 
        \COREAHBLTOAXI_0_AXIMasterIF_RDATA[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(63) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[63]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(62) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[62]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(61) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[61]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(60) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[60]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(59) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[59]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(58) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[58]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(57) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[57]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(56) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[56]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(55) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[55]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(54) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[54]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(53) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[53]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(52) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[52]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(51) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[51]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(50) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[50]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(49) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[49]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(48) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[48]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(47) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[47]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(46) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[46]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(45) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[45]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(44) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[44]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(43) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[43]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(42) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[42]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(41) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[41]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(40) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[40]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(39) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[39]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(38) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[38]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(37) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[37]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(36) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[36]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(35) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[35]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(34) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[34]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(33) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[33]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(32) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[32]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(31) => nc9, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(30) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[30]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(29) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[29]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(28) => nc5, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(27) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[27]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(26) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[26]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(25) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[25]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(24) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[24]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(23) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[23]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(22) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[22]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(21) => nc4, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(20) => nc3, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(19) => nc1, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(18) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[18]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(17) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[17]\, 
        COREAHBLTOAXI_0_AXIMasterIF_WDATA(16) => 
        \COREAHBLTOAXI_0_AXIMasterIF_WDATA[16]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(31) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[31]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(30) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[30]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(29) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[29]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(28) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[28]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(27) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[27]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(26) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[26]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(25) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[25]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(24) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[24]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(23) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[23]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(22) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[22]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(21) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[21]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(20) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[20]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(19) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[19]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(18) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[18]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(17) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[17]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(16) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[16]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(15) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[15]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(14) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[14]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(13) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[13]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(12) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[12]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(11) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[11]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(10) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[10]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(9) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[9]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(8) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[8]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(7) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[7]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(6) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[6]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(5) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[5]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(4) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[4]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(3) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[3]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(2) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[2]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(1) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[1]\, 
        CoreAHBLite_0_AHBmslave10_HWDATA(0) => 
        \CoreAHBLite_0_AHBmslave10_HWDATA[0]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(31) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[31]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(30) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[30]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(29) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[29]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(28) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[28]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(27) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[27]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(26) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[26]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(25) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[25]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(24) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[24]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(23) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[23]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(22) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[22]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(21) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[21]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(20) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[20]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(19) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[19]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(18) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[18]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(17) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[17]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(16) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[16]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(15) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[15]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(14) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[14]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(13) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[13]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(12) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[12]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(11) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[11]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(10) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[10]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(9) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[9]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(8) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[8]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(7) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[7]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(6) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[6]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(5) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[5]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(4) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[4]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(3) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[3]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(2) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[2]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(1) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[1]\, 
        CoreAHBLite_0_AHBmslave10_HRDATA(0) => 
        \CoreAHBLite_0_AHBmslave10_HRDATA[0]\, 
        CoreAHBLite_0_AHBmslave10_HSIZE(1) => 
        \CoreAHBLite_0_AHBmslave10_HSIZE[1]\, 
        CoreAHBLite_0_AHBmslave10_HSIZE(0) => 
        \CoreAHBLite_0_AHBmslave10_HSIZE[0]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(27) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[27]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(26) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[26]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(25) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[25]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(24) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[24]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(23) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[23]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(22) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[22]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(21) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[21]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(20) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[20]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(19) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[19]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(18) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[18]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(17) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[17]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(16) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[16]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(15) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[15]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(14) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[14]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(13) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[13]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(12) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[12]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(11) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[11]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(10) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[10]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(9) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[9]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(8) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[8]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(7) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[7]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(6) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[6]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(5) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[5]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(4) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[4]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(3) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[3]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(2) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[2]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(1) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[1]\, 
        CoreAHBLite_0_AHBmslave10_HADDR(0) => 
        \CoreAHBLite_0_AHBmslave10_HADDR[0]\, 
        COREAHBLTOAXI_0_AXIMasterIF_ARLOCK_0 => 
        \COREAHBLTOAXI_0_AXIMasterIF_ARLOCK[1]\, 
        axi_current_state_0 => \axi_current_state[1]\, 
        axi_current_state_3 => \axi_current_state[4]\, 
        current_state_0 => \current_state[7]\, masterAddrInProg_0
         => \masterAddrInProg[0]\, xhdl1222_0 => \xhdl1222[10]\, 
        MSS_READY => MSS_READY, 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_RREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_WVALID, awaddr_awvalid_clr_d
         => awaddr_awvalid_clr_d, araddr_arvalid_clr_d => 
        araddr_arvalid_clr_d, COREAHBLTOAXI_0_AXIMasterIF_WREADY
         => COREAHBLTOAXI_0_AXIMasterIF_WREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_AWREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_RVALID, 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST => 
        COREAHBLTOAXI_0_AXIMasterIF_RLAST, 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY => 
        COREAHBLTOAXI_0_AXIMasterIF_ARREADY, 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_ARVALID, N_75_i => N_75_i, 
        N_48 => N_48, N_1445_i => N_1445_i, wready_m_xhdl2 => 
        wready_m_xhdl2, N_1446_i => N_1446_i, N_1452_i => 
        N_1452_i, N_1447_i => N_1447_i, N_1451_i => N_1451_i, 
        N_135_i => N_135_i, N_136_i => N_136_i, N_137_i => 
        N_137_i, N_203_i => N_203_i, N_272_i => N_272_i, N_273_i
         => N_273_i, N_274_i => N_274_i, N_275_i => N_275_i, 
        N_276_i => N_276_i, N_277_i => N_277_i, N_382_i => 
        N_382_i, N_381_i => N_381_i, N_278_i => N_278_i, N_380_i
         => N_380_i, N_133_i => N_133_i, N_134_i => N_134_i, 
        N_195_i => N_195_i, N_197_i => N_197_i, N_200_i => 
        N_200_i, N_201_i => N_201_i, N_202_i => N_202_i, N_1450_i
         => N_1450_i, N_1449_i => N_1449_i, N_1448_i => N_1448_i, 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID => 
        COREAHBLTOAXI_0_AXIMasterIF_BVALID, SDRCLK_c => 
        \SDRCLK_c\, CoreAHBLite_0_AHBmslave10_HWRITE => 
        CoreAHBLite_0_AHBmslave10_HWRITE, 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK => 
        CoreAHBLite_0_AHBmslave10_HMASTLOCK, hsel2_0_a2_1 => 
        hsel2_0_a2_1, hsel2 => hsel2, N_91 => N_91, 
        m0PrevDataSlaveReady => m0PrevDataSlaveReady, N_92 => 
        N_92);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity top is

    port( BA           : out   std_logic_vector(1 downto 0);
          CS_N         : out   std_logic_vector(0 to 0);
          DQM          : out   std_logic_vector(1 downto 0);
          SA           : out   std_logic_vector(13 downto 0);
          DQ           : inout std_logic_vector(15 downto 0) := (others => 'Z');
          CAN_RX       : in    std_logic;
          CLK1_PAD     : in    std_logic;
          DEVRST_N     : in    std_logic;
          MMUART_0_RXD : in    std_logic;
          SPI_0_DI     : in    std_logic;
          CAN_TX       : out   std_logic;
          CAN_TX_EN_N  : out   std_logic;
          CAS_N        : out   std_logic;
          CKE          : out   std_logic;
          MMUART_0_TXD : out   std_logic;
          RAS_N        : out   std_logic;
          SDRCLK       : out   std_logic;
          SPI_0_DO     : out   std_logic;
          WE_N         : out   std_logic;
          GPIO_10_BI   : inout std_logic := 'Z';
          GPIO_11_BI   : inout std_logic := 'Z';
          GPIO_12_BI   : inout std_logic := 'Z';
          GPIO_13_BI   : inout std_logic := 'Z';
          GPIO_14_BI   : inout std_logic := 'Z';
          GPIO_15_BI   : inout std_logic := 'Z';
          GPIO_16_BI   : inout std_logic := 'Z';
          GPIO_17_BI   : inout std_logic := 'Z';
          GPIO_18_BI   : inout std_logic := 'Z';
          GPIO_19_BI   : inout std_logic := 'Z';
          GPIO_1_BI    : inout std_logic := 'Z';
          GPIO_20_BI   : inout std_logic := 'Z';
          GPIO_21_BI   : inout std_logic := 'Z';
          GPIO_22_BI   : inout std_logic := 'Z';
          GPIO_23_BI   : inout std_logic := 'Z';
          GPIO_24_BI   : inout std_logic := 'Z';
          GPIO_25_BI   : inout std_logic := 'Z';
          GPIO_26_BI   : inout std_logic := 'Z';
          GPIO_29_BI   : inout std_logic := 'Z';
          GPIO_8_BI    : inout std_logic := 'Z';
          GPIO_9_BI    : inout std_logic := 'Z';
          I2C_0_SCL    : inout std_logic := 'Z';
          I2C_0_SDA    : inout std_logic := 'Z';
          SPI_0_CLK    : inout std_logic := 'Z';
          SPI_0_SS0    : inout std_logic := 'Z'
        );

end top;

architecture DEF_ARCH of top is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component top_sb
    port( DQ_in              : in    std_logic_vector(15 downto 0) := (others => 'U');
          BA_c               : out   std_logic_vector(1 downto 0);
          SA_c               : out   std_logic_vector(11 downto 0);
          sdr_datain_reg     : out   std_logic_vector(15 downto 0);
          DQM_c              : out   std_logic_vector(1 downto 0);
          CS_N_c_0           : out   std_logic;
          CAS_N_c            : out   std_logic;
          CKE_c              : out   std_logic;
          un1_top_sb_0_3_i_i : out   std_logic;
          RAS_N_c            : out   std_logic;
          WE_N_c             : out   std_logic;
          SPI_0_SS0          : inout   std_logic;
          SPI_0_DO           : out   std_logic;
          SPI_0_DI           : in    std_logic := 'U';
          SPI_0_CLK          : inout   std_logic;
          MMUART_0_TXD       : out   std_logic;
          MMUART_0_RXD       : in    std_logic := 'U';
          I2C_0_SDA          : inout   std_logic;
          I2C_0_SCL          : inout   std_logic;
          GPIO_29_BI         : inout   std_logic;
          GPIO_26_BI         : inout   std_logic;
          GPIO_25_BI         : inout   std_logic;
          GPIO_24_BI         : inout   std_logic;
          GPIO_23_BI         : inout   std_logic;
          GPIO_22_BI         : inout   std_logic;
          GPIO_21_BI         : inout   std_logic;
          GPIO_20_BI         : inout   std_logic;
          GPIO_19_BI         : inout   std_logic;
          GPIO_18_BI         : inout   std_logic;
          GPIO_17_BI         : inout   std_logic;
          GPIO_16_BI         : inout   std_logic;
          GPIO_15_BI         : inout   std_logic;
          GPIO_14_BI         : inout   std_logic;
          GPIO_13_BI         : inout   std_logic;
          GPIO_12_BI         : inout   std_logic;
          GPIO_11_BI         : inout   std_logic;
          GPIO_10_BI         : inout   std_logic;
          GPIO_9_BI          : inout   std_logic;
          GPIO_8_BI          : inout   std_logic;
          GPIO_1_BI          : inout   std_logic;
          CAN_TX             : out   std_logic;
          CAN_TX_EN_N        : out   std_logic;
          CAN_RX             : in    std_logic := 'U';
          SDRCLK_c           : out   std_logic;
          CLK1_PAD           : in    std_logic := 'U';
          DEVRST_N           : in    std_logic := 'U'
        );
  end component;

    signal \sdr_datain_reg[0]\, \sdr_datain_reg[1]\, 
        \sdr_datain_reg[2]\, \sdr_datain_reg[3]\, 
        \sdr_datain_reg[4]\, \sdr_datain_reg[5]\, 
        \sdr_datain_reg[6]\, \sdr_datain_reg[7]\, 
        \sdr_datain_reg[8]\, \sdr_datain_reg[9]\, 
        \sdr_datain_reg[10]\, \sdr_datain_reg[11]\, 
        \sdr_datain_reg[12]\, \sdr_datain_reg[13]\, 
        \sdr_datain_reg[14]\, \sdr_datain_reg[15]\, GND_net_1, 
        VCC_net_1, \DQ_in[0]\, \DQ_in[1]\, \DQ_in[2]\, \DQ_in[3]\, 
        \DQ_in[4]\, \DQ_in[5]\, \DQ_in[6]\, \DQ_in[7]\, 
        \DQ_in[8]\, \DQ_in[9]\, \DQ_in[10]\, \DQ_in[11]\, 
        \DQ_in[12]\, \DQ_in[13]\, \DQ_in[14]\, \DQ_in[15]\, 
        \BA_c[0]\, \BA_c[1]\, CAS_N_c, CKE_c, \CS_N_c[0]\, 
        \DQM_c[0]\, \DQM_c[1]\, RAS_N_c, \SA_c[0]\, \SA_c[1]\, 
        \SA_c[2]\, \SA_c[3]\, \SA_c[4]\, \SA_c[5]\, \SA_c[6]\, 
        \SA_c[7]\, \SA_c[8]\, \SA_c[9]\, \SA_c[10]\, \SA_c[11]\, 
        SDRCLK_c, WE_N_c, un1_top_sb_0_3_i_i : std_logic;

    for all : top_sb
	Use entity work.top_sb(DEF_ARCH);
begin 


    WE_N_obuf : OUTBUF
      port map(D => WE_N_c, PAD => WE_N);
    
    \SA_obuf[11]\ : OUTBUF
      port map(D => \SA_c[11]\, PAD => SA(11));
    
    \SA_obuf[13]\ : OUTBUF
      port map(D => GND_net_1, PAD => SA(13));
    
    \DQM_obuf[0]\ : OUTBUF
      port map(D => \DQM_c[0]\, PAD => DQM(0));
    
    \DQ_iobuf[5]\ : BIBUF
      port map(PAD => DQ(5), D => \sdr_datain_reg[5]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[5]\);
    
    \SA_obuf[7]\ : OUTBUF
      port map(D => \SA_c[7]\, PAD => SA(7));
    
    \DQ_iobuf[10]\ : BIBUF
      port map(PAD => DQ(10), D => \sdr_datain_reg[10]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[10]\);
    
    \DQ_iobuf[11]\ : BIBUF
      port map(PAD => DQ(11), D => \sdr_datain_reg[11]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[11]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \DQ_iobuf[0]\ : BIBUF
      port map(PAD => DQ(0), D => \sdr_datain_reg[0]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[0]\);
    
    \SA_obuf[4]\ : OUTBUF
      port map(D => \SA_c[4]\, PAD => SA(4));
    
    \BA_obuf[1]\ : OUTBUF
      port map(D => \BA_c[1]\, PAD => BA(1));
    
    \SA_obuf[3]\ : OUTBUF
      port map(D => \SA_c[3]\, PAD => SA(3));
    
    \DQ_iobuf[1]\ : BIBUF
      port map(PAD => DQ(1), D => \sdr_datain_reg[1]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[1]\);
    
    CKE_obuf : OUTBUF
      port map(D => CKE_c, PAD => CKE);
    
    CAS_N_obuf : OUTBUF
      port map(D => CAS_N_c, PAD => CAS_N);
    
    SDRCLK_obuf : OUTBUF
      port map(D => SDRCLK_c, PAD => SDRCLK);
    
    \DQ_iobuf[14]\ : BIBUF
      port map(PAD => DQ(14), D => \sdr_datain_reg[14]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[14]\);
    
    \SA_obuf[2]\ : OUTBUF
      port map(D => \SA_c[2]\, PAD => SA(2));
    
    \SA_obuf[8]\ : OUTBUF
      port map(D => \SA_c[8]\, PAD => SA(8));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SA_obuf[1]\ : OUTBUF
      port map(D => \SA_c[1]\, PAD => SA(1));
    
    \DQM_obuf[1]\ : OUTBUF
      port map(D => \DQM_c[1]\, PAD => DQM(1));
    
    \DQ_iobuf[8]\ : BIBUF
      port map(PAD => DQ(8), D => \sdr_datain_reg[8]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[8]\);
    
    \DQ_iobuf[13]\ : BIBUF
      port map(PAD => DQ(13), D => \sdr_datain_reg[13]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[13]\);
    
    top_sb_0 : top_sb
      port map(DQ_in(15) => \DQ_in[15]\, DQ_in(14) => \DQ_in[14]\, 
        DQ_in(13) => \DQ_in[13]\, DQ_in(12) => \DQ_in[12]\, 
        DQ_in(11) => \DQ_in[11]\, DQ_in(10) => \DQ_in[10]\, 
        DQ_in(9) => \DQ_in[9]\, DQ_in(8) => \DQ_in[8]\, DQ_in(7)
         => \DQ_in[7]\, DQ_in(6) => \DQ_in[6]\, DQ_in(5) => 
        \DQ_in[5]\, DQ_in(4) => \DQ_in[4]\, DQ_in(3) => 
        \DQ_in[3]\, DQ_in(2) => \DQ_in[2]\, DQ_in(1) => 
        \DQ_in[1]\, DQ_in(0) => \DQ_in[0]\, BA_c(1) => \BA_c[1]\, 
        BA_c(0) => \BA_c[0]\, SA_c(11) => \SA_c[11]\, SA_c(10)
         => \SA_c[10]\, SA_c(9) => \SA_c[9]\, SA_c(8) => 
        \SA_c[8]\, SA_c(7) => \SA_c[7]\, SA_c(6) => \SA_c[6]\, 
        SA_c(5) => \SA_c[5]\, SA_c(4) => \SA_c[4]\, SA_c(3) => 
        \SA_c[3]\, SA_c(2) => \SA_c[2]\, SA_c(1) => \SA_c[1]\, 
        SA_c(0) => \SA_c[0]\, sdr_datain_reg(15) => 
        \sdr_datain_reg[15]\, sdr_datain_reg(14) => 
        \sdr_datain_reg[14]\, sdr_datain_reg(13) => 
        \sdr_datain_reg[13]\, sdr_datain_reg(12) => 
        \sdr_datain_reg[12]\, sdr_datain_reg(11) => 
        \sdr_datain_reg[11]\, sdr_datain_reg(10) => 
        \sdr_datain_reg[10]\, sdr_datain_reg(9) => 
        \sdr_datain_reg[9]\, sdr_datain_reg(8) => 
        \sdr_datain_reg[8]\, sdr_datain_reg(7) => 
        \sdr_datain_reg[7]\, sdr_datain_reg(6) => 
        \sdr_datain_reg[6]\, sdr_datain_reg(5) => 
        \sdr_datain_reg[5]\, sdr_datain_reg(4) => 
        \sdr_datain_reg[4]\, sdr_datain_reg(3) => 
        \sdr_datain_reg[3]\, sdr_datain_reg(2) => 
        \sdr_datain_reg[2]\, sdr_datain_reg(1) => 
        \sdr_datain_reg[1]\, sdr_datain_reg(0) => 
        \sdr_datain_reg[0]\, DQM_c(1) => \DQM_c[1]\, DQM_c(0) => 
        \DQM_c[0]\, CS_N_c_0 => \CS_N_c[0]\, CAS_N_c => CAS_N_c, 
        CKE_c => CKE_c, un1_top_sb_0_3_i_i => un1_top_sb_0_3_i_i, 
        RAS_N_c => RAS_N_c, WE_N_c => WE_N_c, SPI_0_SS0 => 
        SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, 
        SPI_0_CLK => SPI_0_CLK, MMUART_0_TXD => MMUART_0_TXD, 
        MMUART_0_RXD => MMUART_0_RXD, I2C_0_SDA => I2C_0_SDA, 
        I2C_0_SCL => I2C_0_SCL, GPIO_29_BI => GPIO_29_BI, 
        GPIO_26_BI => GPIO_26_BI, GPIO_25_BI => GPIO_25_BI, 
        GPIO_24_BI => GPIO_24_BI, GPIO_23_BI => GPIO_23_BI, 
        GPIO_22_BI => GPIO_22_BI, GPIO_21_BI => GPIO_21_BI, 
        GPIO_20_BI => GPIO_20_BI, GPIO_19_BI => GPIO_19_BI, 
        GPIO_18_BI => GPIO_18_BI, GPIO_17_BI => GPIO_17_BI, 
        GPIO_16_BI => GPIO_16_BI, GPIO_15_BI => GPIO_15_BI, 
        GPIO_14_BI => GPIO_14_BI, GPIO_13_BI => GPIO_13_BI, 
        GPIO_12_BI => GPIO_12_BI, GPIO_11_BI => GPIO_11_BI, 
        GPIO_10_BI => GPIO_10_BI, GPIO_9_BI => GPIO_9_BI, 
        GPIO_8_BI => GPIO_8_BI, GPIO_1_BI => GPIO_1_BI, CAN_TX
         => CAN_TX, CAN_TX_EN_N => CAN_TX_EN_N, CAN_RX => CAN_RX, 
        SDRCLK_c => SDRCLK_c, CLK1_PAD => CLK1_PAD, DEVRST_N => 
        DEVRST_N);
    
    \SA_obuf[5]\ : OUTBUF
      port map(D => \SA_c[5]\, PAD => SA(5));
    
    \DQ_iobuf[9]\ : BIBUF
      port map(PAD => DQ(9), D => \sdr_datain_reg[9]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[9]\);
    
    \DQ_iobuf[3]\ : BIBUF
      port map(PAD => DQ(3), D => \sdr_datain_reg[3]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[3]\);
    
    RAS_N_obuf : OUTBUF
      port map(D => RAS_N_c, PAD => RAS_N);
    
    \SA_obuf[10]\ : OUTBUF
      port map(D => \SA_c[10]\, PAD => SA(10));
    
    \SA_obuf[0]\ : OUTBUF
      port map(D => \SA_c[0]\, PAD => SA(0));
    
    \CS_N_obuf[0]\ : OUTBUF
      port map(D => \CS_N_c[0]\, PAD => CS_N(0));
    
    \BA_obuf[0]\ : OUTBUF
      port map(D => \BA_c[0]\, PAD => BA(0));
    
    \DQ_iobuf[6]\ : BIBUF
      port map(PAD => DQ(6), D => \sdr_datain_reg[6]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[6]\);
    
    \DQ_iobuf[4]\ : BIBUF
      port map(PAD => DQ(4), D => \sdr_datain_reg[4]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[4]\);
    
    \SA_obuf[9]\ : OUTBUF
      port map(D => \SA_c[9]\, PAD => SA(9));
    
    \SA_obuf[6]\ : OUTBUF
      port map(D => \SA_c[6]\, PAD => SA(6));
    
    \DQ_iobuf[15]\ : BIBUF
      port map(PAD => DQ(15), D => \sdr_datain_reg[15]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[15]\);
    
    \DQ_iobuf[7]\ : BIBUF
      port map(PAD => DQ(7), D => \sdr_datain_reg[7]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[7]\);
    
    \DQ_iobuf[2]\ : BIBUF
      port map(PAD => DQ(2), D => \sdr_datain_reg[2]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[2]\);
    
    \DQ_iobuf[12]\ : BIBUF
      port map(PAD => DQ(12), D => \sdr_datain_reg[12]\, E => 
        un1_top_sb_0_3_i_i, Y => \DQ_in[12]\);
    
    \SA_obuf[12]\ : OUTBUF
      port map(D => GND_net_1, PAD => SA(12));
    

end DEF_ARCH; 
